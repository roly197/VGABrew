module font_rom_8x8 (
    input clk,
    input [9:0] addr,
    output reg [7:0] out
);

reg [9:0] addr_r;
always @(posedge clk) begin
  addr_r <= addr;
  case (addr_r)
		10'h000:OUT <=8'b00000000;        
		10'h001:OUT <=8'b00000000;        
		10'h002:OUT <=8'b00000000;        
		10'h003:OUT <=8'b00000000;        
		10'h004:OUT <=8'b00000000;        
		10'h005:OUT <=8'b00000000;        
		10'h006:OUT <=8'b00000000;        
		10'h007:OUT <=8'b00000000;        
		10'h008:OUT <=8'b00000100;        // !
		10'h009:OUT <=8'b00000100;        
		10'h00A:OUT <=8'b00000100;        
		10'h00B:OUT <=8'b00000100;        
		10'h00C:OUT <=8'b00000000;        
		10'h00D:OUT <=8'b00000000;        
		10'h00E:OUT <=8'b00000100;        
		10'h00F:OUT <=8'b00000000;        
		10'h010:OUT <=8'b00001010;        // "
		10'h011:OUT <=8'b00001010;        
		10'h012:OUT <=8'b00001010;        
		10'h013:OUT <=8'b00000000;        
		10'h014:OUT <=8'b00000000;        
		10'h015:OUT <=8'b00000000;        
		10'h016:OUT <=8'b00000000;        
		10'h017:OUT <=8'b00000000;        
		10'h018:OUT <=8'b00001010;        // #
		10'h019:OUT <=8'b00001010;        
		10'h01A:OUT <=8'b00011111;        
		10'h01B:OUT <=8'b00001010;        
		10'h01C:OUT <=8'b00011111;        
		10'h01D:OUT <=8'b00001010;        
		10'h01E:OUT <=8'b00001010;        
		10'h01F:OUT <=8'b00000000;        
		10'h020:OUT <=8'b00000100;        // $
		10'h021:OUT <=8'b00001111;        
		10'h022:OUT <=8'b00010100;        
		10'h023:OUT <=8'b00001110;        
		10'h024:OUT <=8'b00000101;        
		10'h025:OUT <=8'b00011110;        
		10'h026:OUT <=8'b00000100;        
		10'h027:OUT <=8'b00000000;        
		10'h028:OUT <=8'b00011000;        // %
		10'h029:OUT <=8'b00011001;        
		10'h02A:OUT <=8'b00000010;        
		10'h02B:OUT <=8'b00000100;        
		10'h02C:OUT <=8'b00001000;        
		10'h02D:OUT <=8'b00010011;        
		10'h02E:OUT <=8'b00000011;        
		10'h02F:OUT <=8'b00000000;        
		10'h030:OUT <=8'b00001100;        // &
		10'h031:OUT <=8'b00010010;        
		10'h032:OUT <=8'b00010100;        
		10'h033:OUT <=8'b00001000;        
		10'h034:OUT <=8'b00010101;        
		10'h035:OUT <=8'b00010010;        
		10'h036:OUT <=8'b00001101;        
		10'h037:OUT <=8'b00000000;        
		10'h038:OUT <=8'b00001100;        // '
		10'h039:OUT <=8'b00000100;        
		10'h03A:OUT <=8'b00001000;        
		10'h03B:OUT <=8'b00000000;        
		10'h03C:OUT <=8'b00000000;        
		10'h03D:OUT <=8'b00000000;        
		10'h03E:OUT <=8'b00000000;        
		10'h03F:OUT <=8'b00000000;        
		10'h040:OUT <=8'b00000010;        // (
		10'h041:OUT <=8'b00000100;        
		10'h042:OUT <=8'b00001000;        
		10'h043:OUT <=8'b00001000;        
		10'h044:OUT <=8'b00001000;        
		10'h045:OUT <=8'b00000100;        
		10'h046:OUT <=8'b00000010;        
		10'h047:OUT <=8'b00000000;        
		10'h048:OUT <=8'b00001000;        // )
		10'h049:OUT <=8'b00000100;        
		10'h04A:OUT <=8'b00000010;        
		10'h04B:OUT <=8'b00000010;        
		10'h04C:OUT <=8'b00000010;        
		10'h04D:OUT <=8'b00000100;        
		10'h04E:OUT <=8'b00001000;        
		10'h04F:OUT <=8'b00000000;        
		10'h050:OUT <=8'b00000000;        // *
		10'h051:OUT <=8'b00000100;        
		10'h052:OUT <=8'b00010101;        
		10'h053:OUT <=8'b00001110;        
		10'h054:OUT <=8'b00010101;        
		10'h055:OUT <=8'b00000100;        
		10'h056:OUT <=8'b00000000;        
		10'h057:OUT <=8'b00000000;        
		10'h058:OUT <=8'b00000000;        // +
		10'h059:OUT <=8'b00000100;        
		10'h05A:OUT <=8'b00000100;        
		10'h05B:OUT <=8'b00011111;        
		10'h05C:OUT <=8'b00000100;        
		10'h05D:OUT <=8'b00000100;        
		10'h05E:OUT <=8'b00000000;        
		10'h05F:OUT <=8'b00000000;        
		10'h060:OUT <=8'b00000000;        // ,
		10'h061:OUT <=8'b00000000;        
		10'h062:OUT <=8'b00000000;        
		10'h063:OUT <=8'b00000000;        
		10'h064:OUT <=8'b00001100;        
		10'h065:OUT <=8'b00000100;        
		10'h066:OUT <=8'b00001000;        
		10'h067:OUT <=8'b00000000;        
		10'h068:OUT <=8'b00000000;        // -
		10'h069:OUT <=8'b00000000;        
		10'h06A:OUT <=8'b00000000;        
		10'h06B:OUT <=8'b00011111;        
		10'h06C:OUT <=8'b00000000;        
		10'h06D:OUT <=8'b00000000;        
		10'h06E:OUT <=8'b00000000;        
		10'h06F:OUT <=8'b00000000;        
		10'h070:OUT <=8'b00000000;        // .
		10'h071:OUT <=8'b00000000;        
		10'h072:OUT <=8'b00000000;        
		10'h073:OUT <=8'b00000000;        
		10'h074:OUT <=8'b00000000;        
		10'h075:OUT <=8'b00001100;        
		10'h076:OUT <=8'b00001100;        
		10'h077:OUT <=8'b00000000;        
		10'h078:OUT <=8'b00000000;        // /
		10'h079:OUT <=8'b00000001;        
		10'h07A:OUT <=8'b00000010;        
		10'h07B:OUT <=8'b00000100;        
		10'h07C:OUT <=8'b00001000;        
		10'h07D:OUT <=8'b00010000;        
		10'h07E:OUT <=8'b00000000;        
		10'h07F:OUT <=8'b00000000;        
		10'h080:OUT <=8'b00001110;        // 0
		10'h081:OUT <=8'b00010001;        
		10'h082:OUT <=8'b00010011;        
		10'h083:OUT <=8'b00010101;        
		10'h084:OUT <=8'b00011001;        
		10'h085:OUT <=8'b00010001;        
		10'h086:OUT <=8'b00001110;        
		10'h087:OUT <=8'b00000000;        
		10'h088:OUT <=8'b00000100;        // 1
		10'h089:OUT <=8'b00001100;        
		10'h08A:OUT <=8'b00000100;        
		10'h08B:OUT <=8'b00000100;        
		10'h08C:OUT <=8'b00000100;        
		10'h08D:OUT <=8'b00000100;        
		10'h08E:OUT <=8'b00001110;        
		10'h08F:OUT <=8'b00000000;        
		10'h090:OUT <=8'b00001110;        // 2
		10'h091:OUT <=8'b00010001;        
		10'h092:OUT <=8'b00000001;        
		10'h093:OUT <=8'b00000010;        
		10'h094:OUT <=8'b00000100;        
		10'h095:OUT <=8'b00001000;        
		10'h096:OUT <=8'b00011111;        
		10'h097:OUT <=8'b00000000;        
		10'h098:OUT <=8'b00011111;        // 3
		10'h099:OUT <=8'b00000010;        
		10'h09A:OUT <=8'b00000100;        
		10'h09B:OUT <=8'b00000010;        
		10'h09C:OUT <=8'b00000001;        
		10'h09D:OUT <=8'b00010001;        
		10'h09E:OUT <=8'b00001110;        
		10'h09F:OUT <=8'b00000000;        
		10'h0A0:OUT <=8'b00000010;        // 4
		10'h0A1:OUT <=8'b00000110;        
		10'h0A2:OUT <=8'b00001010;        
		10'h0A3:OUT <=8'b00010010;        
		10'h0A4:OUT <=8'b00011111;        
		10'h0A5:OUT <=8'b00000010;        
		10'h0A6:OUT <=8'b00000010;        
		10'h0A7:OUT <=8'b00000000;        
		10'h0A8:OUT <=8'b00011111;        // 5
		10'h0A9:OUT <=8'b00010000;        
		10'h0AA:OUT <=8'b00011110;        
		10'h0AB:OUT <=8'b00000001;        
		10'h0AC:OUT <=8'b00000001;        
		10'h0AD:OUT <=8'b00010001;        
		10'h0AE:OUT <=8'b00001110;        
		10'h0AF:OUT <=8'b00000000;        
		10'h0B0:OUT <=8'b00000110;        // 6
		10'h0B1:OUT <=8'b00001000;        
		10'h0B2:OUT <=8'b00010000;        
		10'h0B3:OUT <=8'b00011110;        
		10'h0B4:OUT <=8'b00010001;        
		10'h0B5:OUT <=8'b00010001;        
		10'h0B6:OUT <=8'b00001110;        
		10'h0B7:OUT <=8'b00000000;        
		10'h0B8:OUT <=8'b00011111;        // 7
		10'h0B9:OUT <=8'b00000001;        
		10'h0BA:OUT <=8'b00000010;        
		10'h0BB:OUT <=8'b00000100;        
		10'h0BC:OUT <=8'b00000100;        
		10'h0BD:OUT <=8'b00000100;        
		10'h0BE:OUT <=8'b00000100;        
		10'h0BF:OUT <=8'b00000000;        
		10'h0C0:OUT <=8'b00011110;        // 8
		10'h0C1:OUT <=8'b00010001;        
		10'h0C2:OUT <=8'b00010001;        
		10'h0C3:OUT <=8'b00001110;        
		10'h0C4:OUT <=8'b00010001;        
		10'h0C5:OUT <=8'b00010001;        
		10'h0C6:OUT <=8'b00001110;        
		10'h0C7:OUT <=8'b00000000;        
		10'h0C8:OUT <=8'b00001110;        // 9
		10'h0C9:OUT <=8'b00010001;        
		10'h0CA:OUT <=8'b00010001;        
		10'h0CB:OUT <=8'b00001111;        
		10'h0CC:OUT <=8'b00000001;        
		10'h0CD:OUT <=8'b00000010;        
		10'h0CE:OUT <=8'b00001100;        
		10'h0CF:OUT <=8'b00000000;        
		10'h0D0:OUT <=8'b00000000;        // :
		10'h0D1:OUT <=8'b00001100;        
		10'h0D2:OUT <=8'b00001100;        
		10'h0D3:OUT <=8'b00000000;        
		10'h0D4:OUT <=8'b00001100;        
		10'h0D5:OUT <=8'b00001100;        
		10'h0D6:OUT <=8'b00000000;        
		10'h0D7:OUT <=8'b00000000;        
		10'h0D8:OUT <=8'b00000000;        // ;
		10'h0D9:OUT <=8'b00001100;        
		10'h0DA:OUT <=8'b00001100;        
		10'h0DB:OUT <=8'b00000000;        
		10'h0DC:OUT <=8'b00001100;        
		10'h0DD:OUT <=8'b00000100;        
		10'h0DE:OUT <=8'b00001000;        
		10'h0DF:OUT <=8'b00000000;        
		10'h0E0:OUT <=8'b00000010;        // <
		10'h0E1:OUT <=8'b00000100;        
		10'h0E2:OUT <=8'b00001000;        
		10'h0E3:OUT <=8'b00010000;        
		10'h0E4:OUT <=8'b00001000;        
		10'h0E5:OUT <=8'b00000100;        
		10'h0E6:OUT <=8'b00000010;        
		10'h0E7:OUT <=8'b00000000;        
		10'h0E8:OUT <=8'b00000000;        // =
		10'h0E9:OUT <=8'b00000000;        
		10'h0EA:OUT <=8'b00011111;        
		10'h0EB:OUT <=8'b00000000;        
		10'h0EC:OUT <=8'b00011111;        
		10'h0ED:OUT <=8'b00000000;        
		10'h0EE:OUT <=8'b00000000;        
		10'h0EF:OUT <=8'b00000000;        
		10'h0F0:OUT <=8'b00001000;        // >
		10'h0F1:OUT <=8'b00000100;        
		10'h0F2:OUT <=8'b00000010;        
		10'h0F3:OUT <=8'b00000001;        
		10'h0F4:OUT <=8'b00000010;        
		10'h0F5:OUT <=8'b00000100;        
		10'h0F6:OUT <=8'b00001000;        
		10'h0F7:OUT <=8'b00000000;        
		10'h0F8:OUT <=8'b00001110;        // ?
		10'h0F9:OUT <=8'b00010001;        
		10'h0FA:OUT <=8'b00000001;        
		10'h0FB:OUT <=8'b00000010;        
		10'h0FC:OUT <=8'b00000100;        
		10'h0FD:OUT <=8'b00000000;        
		10'h0FE:OUT <=8'b00000100;        
		10'h0FF:OUT <=8'b00000000;        
		10'h100:OUT <=8'b00001110;        // @
		10'h101:OUT <=8'b00010001;        
		10'h102:OUT <=8'b00000001;        
		10'h103:OUT <=8'b00001101;        
		10'h104:OUT <=8'b00010101;        
		10'h105:OUT <=8'b00010101;        
		10'h106:OUT <=8'b00001110;        
		10'h107:OUT <=8'b00000000;        
		10'h108:OUT <=8'b00001110;        // A
		10'h109:OUT <=8'b00010001;        
		10'h10A:OUT <=8'b00010001;        
		10'h10B:OUT <=8'b00010001;        
		10'h10C:OUT <=8'b00011111;        
		10'h10D:OUT <=8'b00010001;        
		10'h10E:OUT <=8'b00010001;        
		10'h10F:OUT <=8'b00000000;        
		10'h110:OUT <=8'b00011110;        // B
		10'h111:OUT <=8'b00001001;        
		10'h112:OUT <=8'b00001001;        
		10'h113:OUT <=8'b00001110;        
		10'h114:OUT <=8'b00001001;        
		10'h115:OUT <=8'b00001001;        
		10'h116:OUT <=8'b00011110;        
		10'h117:OUT <=8'b00000000;        
		10'h118:OUT <=8'b00001110;        // C
		10'h119:OUT <=8'b00010001;        
		10'h11A:OUT <=8'b00010000;        
		10'h11B:OUT <=8'b00010000;        
		10'h11C:OUT <=8'b00010000;        
		10'h11D:OUT <=8'b00010001;        
		10'h11E:OUT <=8'b00001110;        
		10'h11F:OUT <=8'b00000000;        
		10'h120:OUT <=8'b00011110;        // D
		10'h121:OUT <=8'b00001001;        
		10'h122:OUT <=8'b00001001;        
		10'h123:OUT <=8'b00001001;        
		10'h124:OUT <=8'b00001001;        
		10'h125:OUT <=8'b00001001;        
		10'h126:OUT <=8'b00011110;        
		10'h127:OUT <=8'b00000000;        
		10'h128:OUT <=8'b00011111;        // E
		10'h129:OUT <=8'b00010000;        
		10'h12A:OUT <=8'b00010000;        
		10'h12B:OUT <=8'b00011111;        
		10'h12C:OUT <=8'b00010000;        
		10'h12D:OUT <=8'b00010000;        
		10'h12E:OUT <=8'b00011111;        
		10'h12F:OUT <=8'b00000000;        
		10'h130:OUT <=8'b00011111;        // F
		10'h131:OUT <=8'b00010000;        
		10'h132:OUT <=8'b00010000;        
		10'h133:OUT <=8'b00011110;        
		10'h134:OUT <=8'b00010000;        
		10'h135:OUT <=8'b00010000;        
		10'h136:OUT <=8'b00010000;        
		10'h137:OUT <=8'b00000000;        
		10'h138:OUT <=8'b00001110;        // G
		10'h139:OUT <=8'b00010001;        
		10'h13A:OUT <=8'b00010000;        
		10'h13B:OUT <=8'b00010011;        
		10'h13C:OUT <=8'b00010001;        
		10'h13D:OUT <=8'b00010001;        
		10'h13E:OUT <=8'b00001111;        
		10'h13F:OUT <=8'b00000000;        
		10'h140:OUT <=8'b00010001;        // H
		10'h141:OUT <=8'b00010001;        
		10'h142:OUT <=8'b00010001;        
		10'h143:OUT <=8'b00011111;        
		10'h144:OUT <=8'b00010001;        
		10'h145:OUT <=8'b00010001;        
		10'h146:OUT <=8'b00010001;        
		10'h147:OUT <=8'b00000000;        
		10'h148:OUT <=8'b00001110;        // I
		10'h149:OUT <=8'b00000100;        
		10'h14A:OUT <=8'b00000100;        
		10'h14B:OUT <=8'b00000100;        
		10'h14C:OUT <=8'b00000100;        
		10'h14D:OUT <=8'b00000100;        
		10'h14E:OUT <=8'b00001110;        
		10'h14F:OUT <=8'b00000000;        
		10'h150:OUT <=8'b00000111;        // J
		10'h151:OUT <=8'b00000010;        
		10'h152:OUT <=8'b00000010;        
		10'h153:OUT <=8'b00000010;        
		10'h154:OUT <=8'b00000010;        
		10'h155:OUT <=8'b00010010;        
		10'h156:OUT <=8'b00001100;        
		10'h157:OUT <=8'b00000000;        
		10'h158:OUT <=8'b00010001;        // K
		10'h159:OUT <=8'b00010010;        
		10'h15A:OUT <=8'b00010100;        
		10'h15B:OUT <=8'b00011000;        
		10'h15C:OUT <=8'b00010100;        
		10'h15D:OUT <=8'b00010010;        
		10'h15E:OUT <=8'b00010001;        
		10'h15F:OUT <=8'b00000000;        
		10'h160:OUT <=8'b00010000;        // L
		10'h161:OUT <=8'b00010000;        
		10'h162:OUT <=8'b00010000;        
		10'h163:OUT <=8'b00010000;        
		10'h164:OUT <=8'b00010000;        
		10'h165:OUT <=8'b00010000;        
		10'h166:OUT <=8'b00011111;        
		10'h167:OUT <=8'b00000000;        
		10'h168:OUT <=8'b00010001;        // M
		10'h169:OUT <=8'b00011011;        
		10'h16A:OUT <=8'b00010101;        
		10'h16B:OUT <=8'b00010101;        
		10'h16C:OUT <=8'b00010001;        
		10'h16D:OUT <=8'b00010001;        
		10'h16E:OUT <=8'b00010001;        
		10'h16F:OUT <=8'b00000000;        
		10'h170:OUT <=8'b00010001;        // N
		10'h171:OUT <=8'b00011001;        
		10'h172:OUT <=8'b00011001;        
		10'h173:OUT <=8'b00010101;        
		10'h174:OUT <=8'b00010011;        
		10'h175:OUT <=8'b00010011;        
		10'h176:OUT <=8'b00010001;        
		10'h177:OUT <=8'b00000000;        
		10'h178:OUT <=8'b00001110;        // O
		10'h179:OUT <=8'b00010001;        
		10'h17A:OUT <=8'b00010001;        
		10'h17B:OUT <=8'b00010001;        
		10'h17C:OUT <=8'b00010001;        
		10'h17D:OUT <=8'b00010001;        
		10'h17E:OUT <=8'b00001110;        
		10'h17F:OUT <=8'b00000000;        
		10'h180:OUT <=8'b00011110;        // P
		10'h181:OUT <=8'b00010001;        
		10'h182:OUT <=8'b00010001;        
		10'h183:OUT <=8'b00011110;        
		10'h184:OUT <=8'b00010000;        
		10'h185:OUT <=8'b00010000;        
		10'h186:OUT <=8'b00010000;        
		10'h187:OUT <=8'b00000000;        
		10'h188:OUT <=8'b00001110;        // Q
		10'h189:OUT <=8'b00010001;        
		10'h18A:OUT <=8'b00010001;        
		10'h18B:OUT <=8'b00010001;        
		10'h18C:OUT <=8'b00010101;        
		10'h18D:OUT <=8'b00010010;        
		10'h18E:OUT <=8'b00011101;        
		10'h18F:OUT <=8'b00000000;        
		10'h190:OUT <=8'b00011110;        // R
		10'h191:OUT <=8'b00010001;        
		10'h192:OUT <=8'b00010001;        
		10'h193:OUT <=8'b00011110;        
		10'h194:OUT <=8'b00010100;        
		10'h195:OUT <=8'b00010010;        
		10'h196:OUT <=8'b00010001;        
		10'h197:OUT <=8'b00000000;        
		10'h198:OUT <=8'b00001110;        // S
		10'h199:OUT <=8'b00010001;        
		10'h19A:OUT <=8'b00010000;        
		10'h19B:OUT <=8'b00001110;        
		10'h19C:OUT <=8'b00000001;        
		10'h19D:OUT <=8'b00010001;        
		10'h19E:OUT <=8'b00001110;        
		10'h19F:OUT <=8'b00000000;        
		10'h1A0:OUT <=8'b00011111;        // T
		10'h1A1:OUT <=8'b00000100;        
		10'h1A2:OUT <=8'b00000100;        
		10'h1A3:OUT <=8'b00000100;        
		10'h1A4:OUT <=8'b00000100;        
		10'h1A5:OUT <=8'b00000100;        
		10'h1A6:OUT <=8'b00000100;        
		10'h1A7:OUT <=8'b00000000;        
		10'h1A8:OUT <=8'b00010001;        // U
		10'h1A9:OUT <=8'b00010001;        
		10'h1AA:OUT <=8'b00010001;        
		10'h1AB:OUT <=8'b00010001;        
		10'h1AC:OUT <=8'b00010001;        
		10'h1AD:OUT <=8'b00010001;        
		10'h1AE:OUT <=8'b00001110;        
		10'h1AF:OUT <=8'b00000000;        
		10'h1B0:OUT <=8'b00010001;        // V
		10'h1B1:OUT <=8'b00010001;        
		10'h1B2:OUT <=8'b00010001;        
		10'h1B3:OUT <=8'b00010001;        
		10'h1B4:OUT <=8'b00010001;        
		10'h1B5:OUT <=8'b00001010;        
		10'h1B6:OUT <=8'b00000100;        
		10'h1B7:OUT <=8'b00000000;        
		10'h1B8:OUT <=8'b00010001;        // W
		10'h1B9:OUT <=8'b00010001;        
		10'h1BA:OUT <=8'b00010001;        
		10'h1BB:OUT <=8'b00010101;        
		10'h1BC:OUT <=8'b00010101;        
		10'h1BD:OUT <=8'b00011011;        
		10'h1BE:OUT <=8'b00010001;        
		10'h1BF:OUT <=8'b00000000;        
		10'h1C0:OUT <=8'b00010001;        // X
		10'h1C1:OUT <=8'b00010001;        
		10'h1C2:OUT <=8'b00001010;        
		10'h1C3:OUT <=8'b00000100;        
		10'h1C4:OUT <=8'b00001010;        
		10'h1C5:OUT <=8'b00010001;        
		10'h1C6:OUT <=8'b00010001;        
		10'h1C7:OUT <=8'b00000000;        
		10'h1C8:OUT <=8'b00010001;        // Y
		10'h1C9:OUT <=8'b00010001;        
		10'h1CA:OUT <=8'b00010001;        
		10'h1CB:OUT <=8'b00001010;        
		10'h1CC:OUT <=8'b00000100;        
		10'h1CD:OUT <=8'b00000100;        
		10'h1CE:OUT <=8'b00000100;        
		10'h1CF:OUT <=8'b00000000;        
		10'h1D0:OUT <=8'b00011111;        // Z
		10'h1D1:OUT <=8'b00000001;        
		10'h1D2:OUT <=8'b00000010;        
		10'h1D3:OUT <=8'b00000100;        
		10'h1D4:OUT <=8'b00001000;        
		10'h1D5:OUT <=8'b00010000;        
		10'h1D6:OUT <=8'b00011111;        
		10'h1D7:OUT <=8'b00000000;        
		10'h1D8:OUT <=8'b00001110;        // [
		10'h1D9:OUT <=8'b00001000;        
		10'h1DA:OUT <=8'b00001000;        
		10'h1DB:OUT <=8'b00001000;        
		10'h1DC:OUT <=8'b00001000;        
		10'h1DD:OUT <=8'b00001000;        
		10'h1DE:OUT <=8'b00001110;        
		10'h1DF:OUT <=8'b00000000;        
		10'h1E0:OUT <=8'b00000000;        // \
		10'h1E1:OUT <=8'b00010000;        
		10'h1E2:OUT <=8'b00001000;        
		10'h1E3:OUT <=8'b00000100;        
		10'h1E4:OUT <=8'b00000010;        
		10'h1E5:OUT <=8'b00000001;        
		10'h1E6:OUT <=8'b00000000;        
		10'h1E7:OUT <=8'b00000000;        
		10'h1E8:OUT <=8'b00001110;        // ]
		10'h1E9:OUT <=8'b00000010;        
		10'h1EA:OUT <=8'b00000010;        
		10'h1EB:OUT <=8'b00000010;        
		10'h1EC:OUT <=8'b00000010;        
		10'h1ED:OUT <=8'b00000010;        
		10'h1EE:OUT <=8'b00001110;        
		10'h1EF:OUT <=8'b00000000;        
		10'h1F0:OUT <=8'b00000100;        // ^
		10'h1F1:OUT <=8'b00001010;        
		10'h1F2:OUT <=8'b00010001;        
		10'h1F3:OUT <=8'b00000000;        
		10'h1F4:OUT <=8'b00000000;        
		10'h1F5:OUT <=8'b00000000;        
		10'h1F6:OUT <=8'b00000000;        
		10'h1F7:OUT <=8'b00000000;        
		10'h1F8:OUT <=8'b00000000;        // _
		10'h1F9:OUT <=8'b00000000;        
		10'h1FA:OUT <=8'b00000000;        
		10'h1FB:OUT <=8'b00000000;        
		10'h1FC:OUT <=8'b00000000;        
		10'h1FD:OUT <=8'b00000000;        
		10'h1FE:OUT <=8'b00011111;        
		10'h1FF:OUT <=8'b00000000;        
		10'h200:OUT <=8'b00010000;        // `
		10'h201:OUT <=8'b00001000;        
		10'h202:OUT <=8'b00000100;        
		10'h203:OUT <=8'b00000000;        
		10'h204:OUT <=8'b00000000;        
		10'h205:OUT <=8'b00000000;        
		10'h206:OUT <=8'b00000000;        
		10'h207:OUT <=8'b00000000;        
		10'h208:OUT <=8'b00000000;        // a
		10'h209:OUT <=8'b00000000;        
		10'h20A:OUT <=8'b00001110;        
		10'h20B:OUT <=8'b00000001;        
		10'h20C:OUT <=8'b00001111;        
		10'h20D:OUT <=8'b00010001;        
		10'h20E:OUT <=8'b00001111;        
		10'h20F:OUT <=8'b00000000;        
		10'h210:OUT <=8'b00010000;        // b
		10'h211:OUT <=8'b00010000;        
		10'h212:OUT <=8'b00010110;        
		10'h213:OUT <=8'b00011001;        
		10'h214:OUT <=8'b00010001;        
		10'h215:OUT <=8'b00010001;        
		10'h216:OUT <=8'b00011110;        
		10'h217:OUT <=8'b00000000;        
		10'h218:OUT <=8'b00000000;        // c
		10'h219:OUT <=8'b00000000;        
		10'h21A:OUT <=8'b00001110;        
		10'h21B:OUT <=8'b00010001;        
		10'h21C:OUT <=8'b00010000;        
		10'h21D:OUT <=8'b00010001;        
		10'h21E:OUT <=8'b00001110;        
		10'h21F:OUT <=8'b00000000;        
		10'h220:OUT <=8'b00000001;        // d
		10'h221:OUT <=8'b00000001;        
		10'h222:OUT <=8'b00001101;        
		10'h223:OUT <=8'b00010011;        
		10'h224:OUT <=8'b00010001;        
		10'h225:OUT <=8'b00010001;        
		10'h226:OUT <=8'b00001111;        
		10'h227:OUT <=8'b00000000;        
		10'h228:OUT <=8'b00000000;        // e
		10'h229:OUT <=8'b00000000;        
		10'h22A:OUT <=8'b00001110;        
		10'h22B:OUT <=8'b00010001;        
		10'h22C:OUT <=8'b00011111;        
		10'h22D:OUT <=8'b00010000;        
		10'h22E:OUT <=8'b00001110;        
		10'h22F:OUT <=8'b00000000;        
		10'h230:OUT <=8'b00000010;        // f
		10'h231:OUT <=8'b00000101;        
		10'h232:OUT <=8'b00000100;        
		10'h233:OUT <=8'b00001110;        
		10'h234:OUT <=8'b00000100;        
		10'h235:OUT <=8'b00000100;        
		10'h236:OUT <=8'b00000100;        
		10'h237:OUT <=8'b00000000;        
		10'h238:OUT <=8'b00000000;        // g
		10'h239:OUT <=8'b00001101;        
		10'h23A:OUT <=8'b00010011;        
		10'h23B:OUT <=8'b00010011;        
		10'h23C:OUT <=8'b00001101;        
		10'h23D:OUT <=8'b00000001;        
		10'h23E:OUT <=8'b00001110;        
		10'h23F:OUT <=8'b00000000;        
		10'h240:OUT <=8'b00010000;        // h
		10'h241:OUT <=8'b00010000;        
		10'h242:OUT <=8'b00010110;        
		10'h243:OUT <=8'b00011001;        
		10'h244:OUT <=8'b00010001;        
		10'h245:OUT <=8'b00010001;        
		10'h246:OUT <=8'b00010001;        
		10'h247:OUT <=8'b00000000;        
		10'h248:OUT <=8'b00000100;        // i
		10'h249:OUT <=8'b00000000;        
		10'h24A:OUT <=8'b00001100;        
		10'h24B:OUT <=8'b00000100;        
		10'h24C:OUT <=8'b00000100;        
		10'h24D:OUT <=8'b00000100;        
		10'h24E:OUT <=8'b00001110;        
		10'h24F:OUT <=8'b00000000;        
		10'h250:OUT <=8'b00000010;        // j
		10'h251:OUT <=8'b00000000;        
		10'h252:OUT <=8'b00000110;        
		10'h253:OUT <=8'b00000010;        
		10'h254:OUT <=8'b00000010;        
		10'h255:OUT <=8'b00010010;        
		10'h256:OUT <=8'b00001100;        
		10'h257:OUT <=8'b00000000;        
		10'h258:OUT <=8'b00001000;        // k
		10'h259:OUT <=8'b00001000;        
		10'h25A:OUT <=8'b00001001;        
		10'h25B:OUT <=8'b00001010;        
		10'h25C:OUT <=8'b00001100;        
		10'h25D:OUT <=8'b00001010;        
		10'h25E:OUT <=8'b00001001;        
		10'h25F:OUT <=8'b00000000;        
		10'h260:OUT <=8'b00001100;        // l
		10'h261:OUT <=8'b00000100;        
		10'h262:OUT <=8'b00000100;        
		10'h263:OUT <=8'b00000100;        
		10'h264:OUT <=8'b00000100;        
		10'h265:OUT <=8'b00000100;        
		10'h266:OUT <=8'b00001110;        
		10'h267:OUT <=8'b00000000;        
		10'h268:OUT <=8'b00000000;        // m
		10'h269:OUT <=8'b00000000;        
		10'h26A:OUT <=8'b00011010;        
		10'h26B:OUT <=8'b00010101;        
		10'h26C:OUT <=8'b00010101;        
		10'h26D:OUT <=8'b00010101;        
		10'h26E:OUT <=8'b00010101;        
		10'h26F:OUT <=8'b00000000;        
		10'h270:OUT <=8'b00000000;        // n
		10'h271:OUT <=8'b00000000;        
		10'h272:OUT <=8'b00010110;        
		10'h273:OUT <=8'b00011001;        
		10'h274:OUT <=8'b00010001;        
		10'h275:OUT <=8'b00010001;        
		10'h276:OUT <=8'b00010001;        
		10'h277:OUT <=8'b00000000;        
		10'h278:OUT <=8'b00000000;        // o
		10'h279:OUT <=8'b00000000;        
		10'h27A:OUT <=8'b00001110;        
		10'h27B:OUT <=8'b00010001;        
		10'h27C:OUT <=8'b00010001;        
		10'h27D:OUT <=8'b00010001;        
		10'h27E:OUT <=8'b00001110;        
		10'h27F:OUT <=8'b00000000;        
		10'h280:OUT <=8'b00000000;        // p
		10'h281:OUT <=8'b00010110;        
		10'h282:OUT <=8'b00011001;        
		10'h283:OUT <=8'b00011001;        
		10'h284:OUT <=8'b00010110;        
		10'h285:OUT <=8'b00010000;        
		10'h286:OUT <=8'b00010000;        
		10'h287:OUT <=8'b00000000;        
		10'h288:OUT <=8'b00000000;        // q
		10'h289:OUT <=8'b00001101;        
		10'h28A:OUT <=8'b00010011;        
		10'h28B:OUT <=8'b00010011;        
		10'h28C:OUT <=8'b00001101;        
		10'h28D:OUT <=8'b00000001;        
		10'h28E:OUT <=8'b00000001;        
		10'h28F:OUT <=8'b00000000;        
		10'h290:OUT <=8'b00000000;        // r
		10'h291:OUT <=8'b00000000;        
		10'h292:OUT <=8'b00010110;        
		10'h293:OUT <=8'b00011001;        
		10'h294:OUT <=8'b00010000;        
		10'h295:OUT <=8'b00010000;        
		10'h296:OUT <=8'b00010000;        
		10'h297:OUT <=8'b00000000;        
		10'h298:OUT <=8'b00000000;        // s
		10'h299:OUT <=8'b00000000;        
		10'h29A:OUT <=8'b00001111;        
		10'h29B:OUT <=8'b00010000;        
		10'h29C:OUT <=8'b00011110;        
		10'h29D:OUT <=8'b00000001;        
		10'h29E:OUT <=8'b00011111;        
		10'h29F:OUT <=8'b00000000;        
		10'h2A0:OUT <=8'b00001000;        // t
		10'h2A1:OUT <=8'b00001000;        
		10'h2A2:OUT <=8'b00011100;        
		10'h2A3:OUT <=8'b00001000;        
		10'h2A4:OUT <=8'b00001000;        
		10'h2A5:OUT <=8'b00001001;        
		10'h2A6:OUT <=8'b00000110;        
		10'h2A7:OUT <=8'b00000000;        
		10'h2A8:OUT <=8'b00000000;        // u
		10'h2A9:OUT <=8'b00000000;        
		10'h2AA:OUT <=8'b00010010;        
		10'h2AB:OUT <=8'b00010010;        
		10'h2AC:OUT <=8'b00010010;        
		10'h2AD:OUT <=8'b00010010;        
		10'h2AE:OUT <=8'b00001101;        
		10'h2AF:OUT <=8'b00000000;        
		10'h2B0:OUT <=8'b00000000;        // v
		10'h2B1:OUT <=8'b00000000;        
		10'h2B2:OUT <=8'b00010001;        
		10'h2B3:OUT <=8'b00010001;        
		10'h2B4:OUT <=8'b00010001;        
		10'h2B5:OUT <=8'b00001010;        
		10'h2B6:OUT <=8'b00000100;        
		10'h2B7:OUT <=8'b00000000;        
		10'h2B8:OUT <=8'b00000000;        // w
		10'h2B9:OUT <=8'b00000000;        
		10'h2BA:OUT <=8'b00010001;        
		10'h2BB:OUT <=8'b00010001;        
		10'h2BC:OUT <=8'b00010101;        
		10'h2BD:OUT <=8'b00010101;        
		10'h2BE:OUT <=8'b00001010;        
		10'h2BF:OUT <=8'b00000000;        
		10'h2C0:OUT <=8'b00000000;        // x
		10'h2C1:OUT <=8'b00000000;        
		10'h2C2:OUT <=8'b00010001;        
		10'h2C3:OUT <=8'b00001010;        
		10'h2C4:OUT <=8'b00000100;        
		10'h2C5:OUT <=8'b00001010;        
		10'h2C6:OUT <=8'b00010001;        
		10'h2C7:OUT <=8'b00000000;        
		10'h2C8:OUT <=8'b00000000;        // y
		10'h2C9:OUT <=8'b00000000;        
		10'h2CA:OUT <=8'b00010001;        
		10'h2CB:OUT <=8'b00010001;        
		10'h2CC:OUT <=8'b00010011;        
		10'h2CD:OUT <=8'b00001101;        
		10'h2CE:OUT <=8'b00000001;        
		10'h2CF:OUT <=8'b00001110;        
		10'h2D0:OUT <=8'b00000000;        // z
		10'h2D1:OUT <=8'b00000000;        
		10'h2D2:OUT <=8'b00011111;        
		10'h2D3:OUT <=8'b00000010;        
		10'h2D4:OUT <=8'b00000100;        
		10'h2D5:OUT <=8'b00001000;        
		10'h2D6:OUT <=8'b00011111;        
		10'h2D7:OUT <=8'b00000000;        
		10'h2D8:OUT <=8'b00000010;        // {
		10'h2D9:OUT <=8'b00000100;        
		10'h2DA:OUT <=8'b00000100;        
		10'h2DB:OUT <=8'b00001000;        
		10'h2DC:OUT <=8'b00000100;        
		10'h2DD:OUT <=8'b00000100;        
		10'h2DE:OUT <=8'b00000010;        
		10'h2DF:OUT <=8'b00000000;        
		10'h2E0:OUT <=8'b00000100;        // |
		10'h2E1:OUT <=8'b00000100;        
		10'h2E2:OUT <=8'b00000100;        
		10'h2E3:OUT <=8'b00000000;        
		10'h2E4:OUT <=8'b00000100;        
		10'h2E5:OUT <=8'b00000100;        
		10'h2E6:OUT <=8'b00000100;        
		10'h2E7:OUT <=8'b00000000;        
		10'h2E8:OUT <=8'b00001000;        // }
		10'h2E9:OUT <=8'b00000100;        
		10'h2EA:OUT <=8'b00000100;        
		10'h2EB:OUT <=8'b00000010;        
		10'h2EC:OUT <=8'b00000100;        
		10'h2ED:OUT <=8'b00000100;        
		10'h2EE:OUT <=8'b00001000;        
		10'h2EF:OUT <=8'b00000000;        
		10'h2F0:OUT <=8'b00001000;        // ~
		10'h2F1:OUT <=8'b00010101;        
		10'h2F2:OUT <=8'b00000010;        
		10'h2F3:OUT <=8'b00000000;        
		10'h2F4:OUT <=8'b00000000;        
		10'h2F5:OUT <=8'b00000000;        
		10'h2F6:OUT <=8'b00000000;        
		10'h2F7:OUT <=8'b00000000;        
    default : out <= 0;
  endcase
end
endmodule
