module font_rom_8x8 (
    input clk,
	 input [6:0] ascii_offset,
	 input [2:0] charpos_y,
    output reg [7:0] out
);

reg [9:0] addr_r;
//assign addr_r = ((ascii_offset << 3) |charpos_y);

always @(posedge clk) begin
  addr_r <= ((ascii_offset << 3) |charpos_y);
  case (addr_r)
		10'h100:out <=8'b00000000;        
		10'h101:out <=8'b00000000;        
		10'h102:out <=8'b00000000;        
		10'h103:out <=8'b00000000;        
		10'h104:out <=8'b00000000;        
		10'h105:out <=8'b00000000;        
		10'h106:out <=8'b00000000;        
		10'h107:out <=8'b00000000;        
		10'h108:out <=8'b00000100;        // !
		10'h109:out <=8'b00000100;        
		10'h10A:out <=8'b00000100;        
		10'h10B:out <=8'b00000100;        
		10'h10C:out <=8'b00000000;        
		10'h10D:out <=8'b00000000;        
		10'h10E:out <=8'b00000100;        
		10'h10F:out <=8'b00000000;        
		10'h110:out <=8'b00001010;        // "
		10'h111:out <=8'b00001010;        
		10'h112:out <=8'b00001010;        
		10'h113:out <=8'b00000000;        
		10'h114:out <=8'b00000000;        
		10'h115:out <=8'b00000000;        
		10'h116:out <=8'b00000000;        
		10'h117:out <=8'b00000000;        
		10'h118:out <=8'b00001010;        // #
		10'h119:out <=8'b00001010;        
		10'h11A:out <=8'b00011111;        
		10'h11B:out <=8'b00001010;        
		10'h11C:out <=8'b00011111;        
		10'h11D:out <=8'b00001010;        
		10'h11E:out <=8'b00001010;        
		10'h11F:out <=8'b00000000;        
		10'h120:out <=8'b00000100;        // $
		10'h121:out <=8'b00001111;        
		10'h122:out <=8'b00010100;        
		10'h123:out <=8'b00001110;        
		10'h124:out <=8'b00000101;        
		10'h125:out <=8'b00011110;        
		10'h126:out <=8'b00000100;        
		10'h127:out <=8'b00000000;        
		10'h128:out <=8'b00011000;        // %
		10'h129:out <=8'b00011001;        
		10'h12A:out <=8'b00000010;        
		10'h12B:out <=8'b00000100;        
		10'h12C:out <=8'b00001000;        
		10'h12D:out <=8'b00010011;        
		10'h12E:out <=8'b00000011;        
		10'h12F:out <=8'b00000000;        
		10'h130:out <=8'b00001100;        // &
		10'h131:out <=8'b00010010;        
		10'h132:out <=8'b00010100;        
		10'h133:out <=8'b00001000;        
		10'h134:out <=8'b00010101;        
		10'h135:out <=8'b00010010;        
		10'h136:out <=8'b00001101;        
		10'h137:out <=8'b00000000;        
		10'h138:out <=8'b00001100;        // '
		10'h139:out <=8'b00000100;        
		10'h13A:out <=8'b00001000;        
		10'h13B:out <=8'b00000000;        
		10'h13C:out <=8'b00000000;        
		10'h13D:out <=8'b00000000;        
		10'h13E:out <=8'b00000000;        
		10'h13F:out <=8'b00000000;        
		10'h140:out <=8'b00000010;        // (
		10'h141:out <=8'b00000100;        
		10'h142:out <=8'b00001000;        
		10'h143:out <=8'b00001000;        
		10'h144:out <=8'b00001000;        
		10'h145:out <=8'b00000100;        
		10'h146:out <=8'b00000010;        
		10'h147:out <=8'b00000000;        
		10'h148:out <=8'b00001000;        // )
		10'h149:out <=8'b00000100;        
		10'h14A:out <=8'b00000010;        
		10'h14B:out <=8'b00000010;        
		10'h14C:out <=8'b00000010;        
		10'h14D:out <=8'b00000100;        
		10'h14E:out <=8'b00001000;        
		10'h14F:out <=8'b00000000;        
		10'h150:out <=8'b00000000;        // *
		10'h151:out <=8'b00000100;        
		10'h152:out <=8'b00010101;        
		10'h153:out <=8'b00001110;        
		10'h154:out <=8'b00010101;        
		10'h155:out <=8'b00000100;        
		10'h156:out <=8'b00000000;        
		10'h157:out <=8'b00000000;        
		10'h158:out <=8'b00000000;        // +
		10'h159:out <=8'b00000100;        
		10'h15A:out <=8'b00000100;        
		10'h15B:out <=8'b00011111;        
		10'h15C:out <=8'b00000100;        
		10'h15D:out <=8'b00000100;        
		10'h15E:out <=8'b00000000;        
		10'h15F:out <=8'b00000000;        
		10'h160:out <=8'b00000000;        // ,
		10'h161:out <=8'b00000000;        
		10'h162:out <=8'b00000000;        
		10'h163:out <=8'b00000000;        
		10'h164:out <=8'b00001100;        
		10'h165:out <=8'b00000100;        
		10'h166:out <=8'b00001000;        
		10'h167:out <=8'b00000000;        
		10'h168:out <=8'b00000000;        // -
		10'h169:out <=8'b00000000;        
		10'h16A:out <=8'b00000000;        
		10'h16B:out <=8'b00011111;        
		10'h16C:out <=8'b00000000;        
		10'h16D:out <=8'b00000000;        
		10'h16E:out <=8'b00000000;        
		10'h16F:out <=8'b00000000;        
		10'h170:out <=8'b00000000;        // .
		10'h171:out <=8'b00000000;        
		10'h172:out <=8'b00000000;        
		10'h173:out <=8'b00000000;        
		10'h174:out <=8'b00000000;        
		10'h175:out <=8'b00001100;        
		10'h176:out <=8'b00001100;        
		10'h177:out <=8'b00000000;        
		10'h178:out <=8'b00000000;        // /
		10'h179:out <=8'b00000001;        
		10'h17A:out <=8'b00000010;        
		10'h17B:out <=8'b00000100;        
		10'h17C:out <=8'b00001000;        
		10'h17D:out <=8'b00010000;        
		10'h17E:out <=8'b00000000;        
		10'h17F:out <=8'b00000000;        
		10'h180:out <=8'b00001110;        // 0
		10'h181:out <=8'b00010001;        
		10'h182:out <=8'b00010011;        
		10'h183:out <=8'b00010101;        
		10'h184:out <=8'b00011001;        
		10'h185:out <=8'b00010001;        
		10'h186:out <=8'b00001110;        
		10'h187:out <=8'b00000000;        
		10'h188:out <=8'b00000100;        // 1
		10'h189:out <=8'b00001100;        
		10'h18A:out <=8'b00000100;        
		10'h18B:out <=8'b00000100;        
		10'h18C:out <=8'b00000100;        
		10'h18D:out <=8'b00000100;        
		10'h18E:out <=8'b00001110;        
		10'h18F:out <=8'b00000000;        
		10'h190:out <=8'b00001110;        // 2
		10'h191:out <=8'b00010001;        
		10'h192:out <=8'b00000001;        
		10'h193:out <=8'b00000010;        
		10'h194:out <=8'b00000100;        
		10'h195:out <=8'b00001000;        
		10'h196:out <=8'b00011111;        
		10'h197:out <=8'b00000000;        
		10'h198:out <=8'b00011111;        // 3
		10'h199:out <=8'b00000010;        
		10'h19A:out <=8'b00000100;        
		10'h19B:out <=8'b00000010;        
		10'h19C:out <=8'b00000001;        
		10'h19D:out <=8'b00010001;        
		10'h19E:out <=8'b00001110;        
		10'h19F:out <=8'b00000000;        
		10'h1A0:out <=8'b00000010;        // 4
		10'h1A1:out <=8'b00000110;        
		10'h1A2:out <=8'b00001010;        
		10'h1A3:out <=8'b00010010;        
		10'h1A4:out <=8'b00011111;        
		10'h1A5:out <=8'b00000010;        
		10'h1A6:out <=8'b00000010;        
		10'h1A7:out <=8'b00000000;        
		10'h1A8:out <=8'b00011111;        // 5
		10'h1A9:out <=8'b00010000;        
		10'h1AA:out <=8'b00011110;        
		10'h1AB:out <=8'b00000001;        
		10'h1AC:out <=8'b00000001;        
		10'h1AD:out <=8'b00010001;        
		10'h1AE:out <=8'b00001110;        
		10'h1AF:out <=8'b00000000;        
		10'h1B0:out <=8'b00000110;        // 6
		10'h1B1:out <=8'b00001000;        
		10'h1B2:out <=8'b00010000;        
		10'h1B3:out <=8'b00011110;        
		10'h1B4:out <=8'b00010001;        
		10'h1B5:out <=8'b00010001;        
		10'h1B6:out <=8'b00001110;        
		10'h1B7:out <=8'b00000000;        
		10'h1B8:out <=8'b00011111;        // 7
		10'h1B9:out <=8'b00000001;        
		10'h1BA:out <=8'b00000010;        
		10'h1BB:out <=8'b00000100;        
		10'h1BC:out <=8'b00000100;        
		10'h1BD:out <=8'b00000100;        
		10'h1BE:out <=8'b00000100;        
		10'h1BF:out <=8'b00000000;        
		10'h1C0:out <=8'b00011110;        // 8
		10'h1C1:out <=8'b00010001;        
		10'h1C2:out <=8'b00010001;        
		10'h1C3:out <=8'b00001110;        
		10'h1C4:out <=8'b00010001;        
		10'h1C5:out <=8'b00010001;        
		10'h1C6:out <=8'b00001110;        
		10'h1C7:out <=8'b00000000;        
		10'h1C8:out <=8'b00001110;        // 9
		10'h1C9:out <=8'b00010001;        
		10'h1CA:out <=8'b00010001;        
		10'h1CB:out <=8'b00001111;        
		10'h1CC:out <=8'b00000001;        
		10'h1CD:out <=8'b00000010;        
		10'h1CE:out <=8'b00001100;        
		10'h1CF:out <=8'b00000000;        
		10'h1D0:out <=8'b00000000;        // :
		10'h1D1:out <=8'b00001100;        
		10'h1D2:out <=8'b00001100;        
		10'h1D3:out <=8'b00000000;        
		10'h1D4:out <=8'b00001100;        
		10'h1D5:out <=8'b00001100;        
		10'h1D6:out <=8'b00000000;        
		10'h1D7:out <=8'b00000000;        
		10'h1D8:out <=8'b00000000;        // ;
		10'h1D9:out <=8'b00001100;        
		10'h1DA:out <=8'b00001100;        
		10'h1DB:out <=8'b00000000;        
		10'h1DC:out <=8'b00001100;        
		10'h1DD:out <=8'b00000100;        
		10'h1DE:out <=8'b00001000;        
		10'h1DF:out <=8'b00000000;        
		10'h1E0:out <=8'b00000010;        // <
		10'h1E1:out <=8'b00000100;        
		10'h1E2:out <=8'b00001000;        
		10'h1E3:out <=8'b00010000;        
		10'h1E4:out <=8'b00001000;        
		10'h1E5:out <=8'b00000100;        
		10'h1E6:out <=8'b00000010;        
		10'h1E7:out <=8'b00000000;        
		10'h1E8:out <=8'b00000000;        // =
		10'h1E9:out <=8'b00000000;        
		10'h1EA:out <=8'b00011111;        
		10'h1EB:out <=8'b00000000;        
		10'h1EC:out <=8'b00011111;        
		10'h1ED:out <=8'b00000000;        
		10'h1EE:out <=8'b00000000;        
		10'h1EF:out <=8'b00000000;        
		10'h1F0:out <=8'b00001000;        // >
		10'h1F1:out <=8'b00000100;        
		10'h1F2:out <=8'b00000010;        
		10'h1F3:out <=8'b00000001;        
		10'h1F4:out <=8'b00000010;        
		10'h1F5:out <=8'b00000100;        
		10'h1F6:out <=8'b00001000;        
		10'h1F7:out <=8'b00000000;        
		10'h1F8:out <=8'b00001110;        // ?
		10'h1F9:out <=8'b00010001;        
		10'h1FA:out <=8'b00000001;        
		10'h1FB:out <=8'b00000010;        
		10'h1FC:out <=8'b00000100;        
		10'h1FD:out <=8'b00000000;        
		10'h1FE:out <=8'b00000100;        
		10'h1FF:out <=8'b00000000;        
		10'h200:out <=8'b00001110;        // @
		10'h201:out <=8'b00010001;        
		10'h202:out <=8'b00000001;        
		10'h203:out <=8'b00001101;        
		10'h204:out <=8'b00010101;        
		10'h205:out <=8'b00010101;        
		10'h206:out <=8'b00001110;        
		10'h207:out <=8'b00000000;        
		10'h208:out <=8'b00001110;        // A
		10'h209:out <=8'b00010001;        
		10'h20A:out <=8'b00010001;        
		10'h20B:out <=8'b00010001;        
		10'h20C:out <=8'b00011111;        
		10'h20D:out <=8'b00010001;        
		10'h20E:out <=8'b00010001;        
		10'h20F:out <=8'b00000000;        
		10'h210:out <=8'b00011110;        // B
		10'h211:out <=8'b00001001;        
		10'h212:out <=8'b00001001;        
		10'h213:out <=8'b00001110;        
		10'h214:out <=8'b00001001;        
		10'h215:out <=8'b00001001;        
		10'h216:out <=8'b00011110;        
		10'h217:out <=8'b00000000;        
		10'h218:out <=8'b00001110;        // C
		10'h219:out <=8'b00010001;        
		10'h21A:out <=8'b00010000;        
		10'h21B:out <=8'b00010000;        
		10'h21C:out <=8'b00010000;        
		10'h21D:out <=8'b00010001;        
		10'h21E:out <=8'b00001110;        
		10'h21F:out <=8'b00000000;        
		10'h220:out <=8'b00011110;        // D
		10'h221:out <=8'b00001001;        
		10'h222:out <=8'b00001001;        
		10'h223:out <=8'b00001001;        
		10'h224:out <=8'b00001001;        
		10'h225:out <=8'b00001001;        
		10'h226:out <=8'b00011110;        
		10'h227:out <=8'b00000000;        
		10'h228:out <=8'b00011111;        // E
		10'h229:out <=8'b00010000;        
		10'h22A:out <=8'b00010000;        
		10'h22B:out <=8'b00011111;        
		10'h22C:out <=8'b00010000;        
		10'h22D:out <=8'b00010000;        
		10'h22E:out <=8'b00011111;        
		10'h22F:out <=8'b00000000;        
		10'h230:out <=8'b00011111;        // F
		10'h231:out <=8'b00010000;        
		10'h232:out <=8'b00010000;        
		10'h233:out <=8'b00011110;        
		10'h234:out <=8'b00010000;        
		10'h235:out <=8'b00010000;        
		10'h236:out <=8'b00010000;        
		10'h237:out <=8'b00000000;        
		10'h238:out <=8'b00001110;        // G
		10'h239:out <=8'b00010001;        
		10'h23A:out <=8'b00010000;        
		10'h23B:out <=8'b00010011;        
		10'h23C:out <=8'b00010001;        
		10'h23D:out <=8'b00010001;        
		10'h23E:out <=8'b00001111;        
		10'h23F:out <=8'b00000000;        
		10'h240:out <=8'b00010001;        // H
		10'h241:out <=8'b00010001;        
		10'h242:out <=8'b00010001;        
		10'h243:out <=8'b00011111;        
		10'h244:out <=8'b00010001;        
		10'h245:out <=8'b00010001;        
		10'h246:out <=8'b00010001;        
		10'h247:out <=8'b00000000;        
		10'h248:out <=8'b00001110;        // I
		10'h249:out <=8'b00000100;        
		10'h24A:out <=8'b00000100;        
		10'h24B:out <=8'b00000100;        
		10'h24C:out <=8'b00000100;        
		10'h24D:out <=8'b00000100;        
		10'h24E:out <=8'b00001110;        
		10'h24F:out <=8'b00000000;        
		10'h250:out <=8'b00000111;        // J
		10'h251:out <=8'b00000010;        
		10'h252:out <=8'b00000010;        
		10'h253:out <=8'b00000010;        
		10'h254:out <=8'b00000010;        
		10'h255:out <=8'b00010010;        
		10'h256:out <=8'b00001100;        
		10'h257:out <=8'b00000000;        
		10'h258:out <=8'b00010001;        // K
		10'h259:out <=8'b00010010;        
		10'h25A:out <=8'b00010100;        
		10'h25B:out <=8'b00011000;        
		10'h25C:out <=8'b00010100;        
		10'h25D:out <=8'b00010010;        
		10'h25E:out <=8'b00010001;        
		10'h25F:out <=8'b00000000;        
		10'h260:out <=8'b00010000;        // L
		10'h261:out <=8'b00010000;        
		10'h262:out <=8'b00010000;        
		10'h263:out <=8'b00010000;        
		10'h264:out <=8'b00010000;        
		10'h265:out <=8'b00010000;        
		10'h266:out <=8'b00011111;        
		10'h267:out <=8'b00000000;        
		10'h268:out <=8'b00010001;        // M
		10'h269:out <=8'b00011011;        
		10'h26A:out <=8'b00010101;        
		10'h26B:out <=8'b00010101;        
		10'h26C:out <=8'b00010001;        
		10'h26D:out <=8'b00010001;        
		10'h26E:out <=8'b00010001;        
		10'h26F:out <=8'b00000000;        
		10'h270:out <=8'b00010001;        // N
		10'h271:out <=8'b00011001;        
		10'h272:out <=8'b00011001;        
		10'h273:out <=8'b00010101;        
		10'h274:out <=8'b00010011;        
		10'h275:out <=8'b00010011;        
		10'h276:out <=8'b00010001;        
		10'h277:out <=8'b00000000;        
		10'h278:out <=8'b00001110;        // O
		10'h279:out <=8'b00010001;        
		10'h27A:out <=8'b00010001;        
		10'h27B:out <=8'b00010001;        
		10'h27C:out <=8'b00010001;        
		10'h27D:out <=8'b00010001;        
		10'h27E:out <=8'b00001110;        
		10'h27F:out <=8'b00000000;        
		10'h280:out <=8'b00011110;        // P
		10'h281:out <=8'b00010001;        
		10'h282:out <=8'b00010001;        
		10'h283:out <=8'b00011110;        
		10'h284:out <=8'b00010000;        
		10'h285:out <=8'b00010000;        
		10'h286:out <=8'b00010000;        
		10'h287:out <=8'b00000000;        
		10'h288:out <=8'b00001110;        // Q
		10'h289:out <=8'b00010001;        
		10'h28A:out <=8'b00010001;        
		10'h28B:out <=8'b00010001;        
		10'h28C:out <=8'b00010101;        
		10'h28D:out <=8'b00010010;        
		10'h28E:out <=8'b00011101;        
		10'h28F:out <=8'b00000000;        
		10'h290:out <=8'b00011110;        // R
		10'h291:out <=8'b00010001;        
		10'h292:out <=8'b00010001;        
		10'h293:out <=8'b00011110;        
		10'h294:out <=8'b00010100;        
		10'h295:out <=8'b00010010;        
		10'h296:out <=8'b00010001;        
		10'h297:out <=8'b00000000;        
		10'h298:out <=8'b00001110;        // S
		10'h299:out <=8'b00010001;        
		10'h29A:out <=8'b00010000;        
		10'h29B:out <=8'b00001110;        
		10'h29C:out <=8'b00000001;        
		10'h29D:out <=8'b00010001;        
		10'h29E:out <=8'b00001110;        
		10'h29F:out <=8'b00000000;        
		10'h2A0:out <=8'b00011111;        // T
		10'h2A1:out <=8'b00000100;        
		10'h2A2:out <=8'b00000100;        
		10'h2A3:out <=8'b00000100;        
		10'h2A4:out <=8'b00000100;        
		10'h2A5:out <=8'b00000100;        
		10'h2A6:out <=8'b00000100;        
		10'h2A7:out <=8'b00000000;        
		10'h2A8:out <=8'b00010001;        // U
		10'h2A9:out <=8'b00010001;        
		10'h2AA:out <=8'b00010001;        
		10'h2AB:out <=8'b00010001;        
		10'h2AC:out <=8'b00010001;        
		10'h2AD:out <=8'b00010001;        
		10'h2AE:out <=8'b00001110;        
		10'h2AF:out <=8'b00000000;        
		10'h2B0:out <=8'b00010001;        // V
		10'h2B1:out <=8'b00010001;        
		10'h2B2:out <=8'b00010001;        
		10'h2B3:out <=8'b00010001;        
		10'h2B4:out <=8'b00010001;        
		10'h2B5:out <=8'b00001010;        
		10'h2B6:out <=8'b00000100;        
		10'h2B7:out <=8'b00000000;        
		10'h2B8:out <=8'b00010001;        // W
		10'h2B9:out <=8'b00010001;        
		10'h2BA:out <=8'b00010001;        
		10'h2BB:out <=8'b00010101;        
		10'h2BC:out <=8'b00010101;        
		10'h2BD:out <=8'b00011011;        
		10'h2BE:out <=8'b00010001;        
		10'h2BF:out <=8'b00000000;        
		10'h2C0:out <=8'b00010001;        // X
		10'h2C1:out <=8'b00010001;        
		10'h2C2:out <=8'b00001010;        
		10'h2C3:out <=8'b00000100;        
		10'h2C4:out <=8'b00001010;        
		10'h2C5:out <=8'b00010001;        
		10'h2C6:out <=8'b00010001;        
		10'h2C7:out <=8'b00000000;        
		10'h2C8:out <=8'b00010001;        // Y
		10'h2C9:out <=8'b00010001;        
		10'h2CA:out <=8'b00010001;        
		10'h2CB:out <=8'b00001010;        
		10'h2CC:out <=8'b00000100;        
		10'h2CD:out <=8'b00000100;        
		10'h2CE:out <=8'b00000100;        
		10'h2CF:out <=8'b00000000;        
		10'h2D0:out <=8'b00011111;        // Z
		10'h2D1:out <=8'b00000001;        
		10'h2D2:out <=8'b00000010;        
		10'h2D3:out <=8'b00000100;        
		10'h2D4:out <=8'b00001000;        
		10'h2D5:out <=8'b00010000;        
		10'h2D6:out <=8'b00011111;        
		10'h2D7:out <=8'b00000000;        
		10'h2D8:out <=8'b00001110;        // [
		10'h2D9:out <=8'b00001000;        
		10'h2DA:out <=8'b00001000;        
		10'h2DB:out <=8'b00001000;        
		10'h2DC:out <=8'b00001000;        
		10'h2DD:out <=8'b00001000;        
		10'h2DE:out <=8'b00001110;        
		10'h2DF:out <=8'b00000000;        
		10'h2E0:out <=8'b00000000;        // \
		10'h2E1:out <=8'b00010000;        
		10'h2E2:out <=8'b00001000;        
		10'h2E3:out <=8'b00000100;        
		10'h2E4:out <=8'b00000010;        
		10'h2E5:out <=8'b00000001;        
		10'h2E6:out <=8'b00000000;        
		10'h2E7:out <=8'b00000000;        
		10'h2E8:out <=8'b00001110;        // ]
		10'h2E9:out <=8'b00000010;        
		10'h2EA:out <=8'b00000010;        
		10'h2EB:out <=8'b00000010;        
		10'h2EC:out <=8'b00000010;        
		10'h2ED:out <=8'b00000010;        
		10'h2EE:out <=8'b00001110;        
		10'h2EF:out <=8'b00000000;        
		10'h2F0:out <=8'b00000100;        // ^
		10'h2F1:out <=8'b00001010;        
		10'h2F2:out <=8'b00010001;        
		10'h2F3:out <=8'b00000000;        
		10'h2F4:out <=8'b00000000;        
		10'h2F5:out <=8'b00000000;        
		10'h2F6:out <=8'b00000000;        
		10'h2F7:out <=8'b00000000;        
		10'h2F8:out <=8'b00000000;        // _
		10'h2F9:out <=8'b00000000;        
		10'h2FA:out <=8'b00000000;        
		10'h2FB:out <=8'b00000000;        
		10'h2FC:out <=8'b00000000;        
		10'h2FD:out <=8'b00000000;        
		10'h2FE:out <=8'b00011111;        
		10'h2FF:out <=8'b00000000;        
		10'h300:out <=8'b00010000;        // `
		10'h301:out <=8'b00001000;        
		10'h302:out <=8'b00000100;        
		10'h303:out <=8'b00000000;        
		10'h304:out <=8'b00000000;        
		10'h305:out <=8'b00000000;        
		10'h306:out <=8'b00000000;        
		10'h307:out <=8'b00000000;        
		10'h308:out <=8'b00000000;        // a
		10'h309:out <=8'b00000000;        
		10'h30A:out <=8'b00001110;        
		10'h30B:out <=8'b00000001;        
		10'h30C:out <=8'b00001111;        
		10'h30D:out <=8'b00010001;        
		10'h30E:out <=8'b00001111;        
		10'h30F:out <=8'b00000000;        
		10'h310:out <=8'b00010000;        // b
		10'h311:out <=8'b00010000;        
		10'h312:out <=8'b00010110;        
		10'h313:out <=8'b00011001;        
		10'h314:out <=8'b00010001;        
		10'h315:out <=8'b00010001;        
		10'h316:out <=8'b00011110;        
		10'h317:out <=8'b00000000;        
		10'h318:out <=8'b00000000;        // c
		10'h319:out <=8'b00000000;        
		10'h31A:out <=8'b00001110;        
		10'h31B:out <=8'b00010001;        
		10'h31C:out <=8'b00010000;        
		10'h31D:out <=8'b00010001;        
		10'h31E:out <=8'b00001110;        
		10'h31F:out <=8'b00000000;        
		10'h320:out <=8'b00000001;        // d
		10'h321:out <=8'b00000001;        
		10'h322:out <=8'b00001101;        
		10'h323:out <=8'b00010011;        
		10'h324:out <=8'b00010001;        
		10'h325:out <=8'b00010001;        
		10'h326:out <=8'b00001111;        
		10'h327:out <=8'b00000000;        
		10'h328:out <=8'b00000000;        // e
		10'h329:out <=8'b00000000;        
		10'h32A:out <=8'b00001110;        
		10'h32B:out <=8'b00010001;        
		10'h32C:out <=8'b00011111;        
		10'h32D:out <=8'b00010000;        
		10'h32E:out <=8'b00001110;        
		10'h32F:out <=8'b00000000;        
		10'h330:out <=8'b00000010;        // f
		10'h331:out <=8'b00000101;        
		10'h332:out <=8'b00000100;        
		10'h333:out <=8'b00001110;        
		10'h334:out <=8'b00000100;        
		10'h335:out <=8'b00000100;        
		10'h336:out <=8'b00000100;        
		10'h337:out <=8'b00000000;        
		10'h338:out <=8'b00000000;        // g
		10'h339:out <=8'b00001101;        
		10'h33A:out <=8'b00010011;        
		10'h33B:out <=8'b00010011;        
		10'h33C:out <=8'b00001101;        
		10'h33D:out <=8'b00000001;        
		10'h33E:out <=8'b00001110;        
		10'h33F:out <=8'b00000000;        
		10'h340:out <=8'b00010000;        // h
		10'h341:out <=8'b00010000;        
		10'h342:out <=8'b00010110;        
		10'h343:out <=8'b00011001;        
		10'h344:out <=8'b00010001;        
		10'h345:out <=8'b00010001;        
		10'h346:out <=8'b00010001;        
		10'h347:out <=8'b00000000;        
		10'h348:out <=8'b00000100;        // i
		10'h349:out <=8'b00000000;        
		10'h34A:out <=8'b00001100;        
		10'h34B:out <=8'b00000100;        
		10'h34C:out <=8'b00000100;        
		10'h34D:out <=8'b00000100;        
		10'h34E:out <=8'b00001110;        
		10'h34F:out <=8'b00000000;        
		10'h350:out <=8'b00000010;        // j
		10'h351:out <=8'b00000000;        
		10'h352:out <=8'b00000110;        
		10'h353:out <=8'b00000010;        
		10'h354:out <=8'b00000010;        
		10'h355:out <=8'b00010010;        
		10'h356:out <=8'b00001100;        
		10'h357:out <=8'b00000000;        
		10'h358:out <=8'b00001000;        // k
		10'h359:out <=8'b00001000;        
		10'h35A:out <=8'b00001001;        
		10'h35B:out <=8'b00001010;        
		10'h35C:out <=8'b00001100;        
		10'h35D:out <=8'b00001010;        
		10'h35E:out <=8'b00001001;        
		10'h35F:out <=8'b00000000;        
		10'h360:out <=8'b00001100;        // l
		10'h361:out <=8'b00000100;        
		10'h362:out <=8'b00000100;        
		10'h363:out <=8'b00000100;        
		10'h364:out <=8'b00000100;        
		10'h365:out <=8'b00000100;        
		10'h366:out <=8'b00001110;        
		10'h367:out <=8'b00000000;        
		10'h368:out <=8'b00000000;        // m
		10'h369:out <=8'b00000000;        
		10'h36A:out <=8'b00011010;        
		10'h36B:out <=8'b00010101;        
		10'h36C:out <=8'b00010101;        
		10'h36D:out <=8'b00010101;        
		10'h36E:out <=8'b00010101;        
		10'h36F:out <=8'b00000000;        
		10'h370:out <=8'b00000000;        // n
		10'h371:out <=8'b00000000;        
		10'h372:out <=8'b00010110;        
		10'h373:out <=8'b00011001;        
		10'h374:out <=8'b00010001;        
		10'h375:out <=8'b00010001;        
		10'h376:out <=8'b00010001;        
		10'h377:out <=8'b00000000;        
		10'h378:out <=8'b00000000;        // o
		10'h379:out <=8'b00000000;        
		10'h37A:out <=8'b00001110;        
		10'h37B:out <=8'b00010001;        
		10'h37C:out <=8'b00010001;        
		10'h37D:out <=8'b00010001;        
		10'h37E:out <=8'b00001110;        
		10'h37F:out <=8'b00000000;        
		10'h380:out <=8'b00000000;        // p
		10'h381:out <=8'b00010110;        
		10'h382:out <=8'b00011001;        
		10'h383:out <=8'b00011001;        
		10'h384:out <=8'b00010110;        
		10'h385:out <=8'b00010000;        
		10'h386:out <=8'b00010000;        
		10'h387:out <=8'b00000000;        
		10'h388:out <=8'b00000000;        // q
		10'h389:out <=8'b00001101;        
		10'h38A:out <=8'b00010011;        
		10'h38B:out <=8'b00010011;        
		10'h38C:out <=8'b00001101;        
		10'h38D:out <=8'b00000001;        
		10'h38E:out <=8'b00000001;        
		10'h38F:out <=8'b00000000;        
		10'h390:out <=8'b00000000;        // r
		10'h391:out <=8'b00000000;        
		10'h392:out <=8'b00010110;        
		10'h393:out <=8'b00011001;        
		10'h394:out <=8'b00010000;        
		10'h395:out <=8'b00010000;        
		10'h396:out <=8'b00010000;        
		10'h397:out <=8'b00000000;        
		10'h398:out <=8'b00000000;        // s
		10'h399:out <=8'b00000000;        
		10'h39A:out <=8'b00001111;        
		10'h39B:out <=8'b00010000;        
		10'h39C:out <=8'b00011110;        
		10'h39D:out <=8'b00000001;        
		10'h39E:out <=8'b00011111;        
		10'h39F:out <=8'b00000000;        
		10'h3A0:out <=8'b00001000;        // t
		10'h3A1:out <=8'b00001000;        
		10'h3A2:out <=8'b00011100;        
		10'h3A3:out <=8'b00001000;        
		10'h3A4:out <=8'b00001000;        
		10'h3A5:out <=8'b00001001;        
		10'h3A6:out <=8'b00000110;        
		10'h3A7:out <=8'b00000000;        
		10'h3A8:out <=8'b00000000;        // u
		10'h3A9:out <=8'b00000000;        
		10'h3AA:out <=8'b00010010;        
		10'h3AB:out <=8'b00010010;        
		10'h3AC:out <=8'b00010010;        
		10'h3AD:out <=8'b00010010;        
		10'h3AE:out <=8'b00001101;        
		10'h3AF:out <=8'b00000000;        
		10'h3B0:out <=8'b00000000;        // v
		10'h3B1:out <=8'b00000000;        
		10'h3B2:out <=8'b00010001;        
		10'h3B3:out <=8'b00010001;        
		10'h3B4:out <=8'b00010001;        
		10'h3B5:out <=8'b00001010;        
		10'h3B6:out <=8'b00000100;        
		10'h3B7:out <=8'b00000000;        
		10'h3B8:out <=8'b00000000;        // w
		10'h3B9:out <=8'b00000000;        
		10'h3BA:out <=8'b00010001;        
		10'h3BB:out <=8'b00010001;        
		10'h3BC:out <=8'b00010101;        
		10'h3BD:out <=8'b00010101;        
		10'h3BE:out <=8'b00001010;        
		10'h3BF:out <=8'b00000000;        
		10'h3C0:out <=8'b00000000;        // x
		10'h3C1:out <=8'b00000000;        
		10'h3C2:out <=8'b00010001;        
		10'h3C3:out <=8'b00001010;        
		10'h3C4:out <=8'b00000100;        
		10'h3C5:out <=8'b00001010;        
		10'h3C6:out <=8'b00010001;        
		10'h3C7:out <=8'b00000000;        
		10'h3C8:out <=8'b00000000;        // y
		10'h3C9:out <=8'b00000000;        
		10'h3CA:out <=8'b00010001;        
		10'h3CB:out <=8'b00010001;        
		10'h3CC:out <=8'b00010011;        
		10'h3CD:out <=8'b00001101;        
		10'h3CE:out <=8'b00000001;        
		10'h3CF:out <=8'b00001110;        
		10'h3D0:out <=8'b00000000;        // z
		10'h3D1:out <=8'b00000000;        
		10'h3D2:out <=8'b00011111;        
		10'h3D3:out <=8'b00000010;        
		10'h3D4:out <=8'b00000100;        
		10'h3D5:out <=8'b00001000;        
		10'h3D6:out <=8'b00011111;        
		10'h3D7:out <=8'b00000000;        
		10'h3D8:out <=8'b00000010;        // {
		10'h3D9:out <=8'b00000100;        
		10'h3DA:out <=8'b00000100;        
		10'h3DB:out <=8'b00001000;        
		10'h3DC:out <=8'b00000100;        
		10'h3DD:out <=8'b00000100;        
		10'h3DE:out <=8'b00000010;        
		10'h3DF:out <=8'b00000000;        
		10'h3E0:out <=8'b00000100;        // |
		10'h3E1:out <=8'b00000100;        
		10'h3E2:out <=8'b00000100;        
		10'h3E3:out <=8'b00000000;        
		10'h3E4:out <=8'b00000100;        
		10'h3E5:out <=8'b00000100;        
		10'h3E6:out <=8'b00000100;        
		10'h3E7:out <=8'b00000000;        
		10'h3E8:out <=8'b00001000;        // }
		10'h3E9:out <=8'b00000100;        
		10'h3EA:out <=8'b00000100;        
		10'h3EB:out <=8'b00000010;        
		10'h3EC:out <=8'b00000100;        
		10'h3ED:out <=8'b00000100;        
		10'h3EE:out <=8'b00001000;        
		10'h3EF:out <=8'b00000000;        
		10'h3F0:out <=8'b00001000;        // ~
		10'h3F1:out <=8'b00010101;        
		10'h3F2:out <=8'b00000010;        
		10'h3F3:out <=8'b00000000;        
		10'h3F4:out <=8'b00000000;        
		10'h3F5:out <=8'b00000000;        
		10'h3F6:out <=8'b00000000;        
		10'h3F7:out <=8'b00000000;               
    default : out <= 0;
  endcase
end
endmodule
