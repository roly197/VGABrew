module font_rom_8x8 (
    input clk,
	 input [6:0] ascii_offset,
	 input [2:0] charpos_y,
    output reg [7:0] out
);

reg [9:0] addr_r;
//assign addr_r = ((ascii_offset << 3) |charpos_y);

always @(posedge clk) begin
  addr_r <= ((ascii_offset << 3) |charpos_y);
  case (addr_r)
		10'h100:out <=8'b00000000;        
		10'h101:out <=8'b00000000;        
		10'h102:out <=8'b00000000;        
		10'h103:out <=8'b00000000;        
		10'h104:out <=8'b00000000;        
		10'h105:out <=8'b00000000;        
		10'h106:out <=8'b00000000;        
		10'h107:out <=8'b00000000;        
		10'h108:out <=8'b00000100;        // !
		10'h109:out <=8'b00000100;        
		10'h10A:out <=8'b00000100;        
		10'h10B:out <=8'b00000100;        
		10'h10C:out <=8'b00000000;        
		10'h10D:out <=8'b00000000;        
		10'h10E:out <=8'b00000100;        
		10'h10F:out <=8'b00000000;        
		10'h110:out <=8'b00001010;        // "
		10'h111:out <=8'b00001010;        
		10'h112:out <=8'b00001010;        
		10'h113:out <=8'b00000000;        
		10'h114:out <=8'b00000000;        
		10'h115:out <=8'b00000000;        
		10'h116:out <=8'b00000000;        
		10'h117:out <=8'b00000000;        
		10'h118:out <=8'b00001010;        // #
		10'h119:out <=8'b00001010;        
		10'h11A:out <=8'b00011111;        
		10'h11B:out <=8'b00001010;        
		10'h11C:out <=8'b00011111;        
		10'h11D:out <=8'b00001010;        
		10'h11E:out <=8'b00001010;        
		10'h11F:out <=8'b00000000;        
		10'h120:out <=8'b00000100;        // $
		10'h121:out <=8'b00001111;        
		10'h122:out <=8'b00010100;        
		10'h123:out <=8'b00001110;        
		10'h124:out <=8'b00000101;        
		10'h125:out <=8'b00011110;        
		10'h126:out <=8'b00000100;        
		10'h127:out <=8'b00000000;        
		10'h128:out <=8'b00011000;        // %
		10'h129:out <=8'b00011001;        
		10'h12A:out <=8'b00000010;        
		10'h12B:out <=8'b00000100;        
		10'h12C:out <=8'b00001000;        
		10'h12D:out <=8'b00010011;        
		10'h12E:out <=8'b00000011;        
		10'h12F:out <=8'b00000000;        
		10'h130:out <=8'b00001100;        // &
		10'h131:out <=8'b00010010;        
		10'h132:out <=8'b00010100;        
		10'h133:out <=8'b00001000;        
		10'h134:out <=8'b00010101;        
		10'h135:out <=8'b00010010;        
		10'h136:out <=8'b00001101;        
		10'h137:out <=8'b00000000;        
		10'h138:out <=8'b00001100;        // '
		10'h139:out <=8'b00000100;        
		10'h13A:out <=8'b00001000;        
		10'h13B:out <=8'b00000000;        
		10'h13C:out <=8'b00000000;        
		10'h13D:out <=8'b00000000;        
		10'h13E:out <=8'b00000000;        
		10'h13F:out <=8'b00000000;        
		10'h140:out <=8'b00000010;        // (
		10'h141:out <=8'b00000100;        
		10'h142:out <=8'b00001000;        
		10'h143:out <=8'b00001000;        
		10'h144:out <=8'b00001000;        
		10'h145:out <=8'b00000100;        
		10'h146:out <=8'b00000010;        
		10'h147:out <=8'b00000000;        
		10'h148:out <=8'b00001000;        // )
		10'h149:out <=8'b00000100;        
		10'h14A:out <=8'b00000010;        
		10'h14B:out <=8'b00000010;        
		10'h14C:out <=8'b00000010;        
		10'h14D:out <=8'b00000100;        
		10'h14E:out <=8'b00001000;        
		10'h14F:out <=8'b00000000;        
		10'h150:out <=8'b00000000;        // *
		10'h151:out <=8'b00000100;        
		10'h152:out <=8'b00010101;        
		10'h153:out <=8'b00001110;        
		10'h154:out <=8'b00010101;        
		10'h155:out <=8'b00000100;        
		10'h156:out <=8'b00000000;        
		10'h157:out <=8'b00000000;        
		10'h158:out <=8'b00000000;        // +
		10'h159:out <=8'b00000100;        
		10'h15A:out <=8'b00000100;        
		10'h15B:out <=8'b00011111;        
		10'h15C:out <=8'b00000100;        
		10'h15D:out <=8'b00000100;        
		10'h15E:out <=8'b00000000;        
		10'h15F:out <=8'b00000000;        
		10'h160:out <=8'b00000000;        // ,
		10'h161:out <=8'b00000000;        
		10'h162:out <=8'b00000000;        
		10'h163:out <=8'b00000000;        
		10'h164:out <=8'b00001100;        
		10'h165:out <=8'b00000100;        
		10'h166:out <=8'b00001000;        
		10'h167:out <=8'b00000000;        
		10'h168:out <=8'b00000000;        // -
		10'h169:out <=8'b00000000;        
		10'h16A:out <=8'b00000000;        
		10'h16B:out <=8'b00011111;        
		10'h16C:out <=8'b00000000;        
		10'h16D:out <=8'b00000000;        
		10'h16E:out <=8'b00000000;        
		10'h16F:out <=8'b00000000;        
		10'h170:out <=8'b00000000;        // .
		10'h171:out <=8'b00000000;        
		10'h172:out <=8'b00000000;        
		10'h173:out <=8'b00000000;        
		10'h174:out <=8'b00000000;        
		10'h175:out <=8'b00001100;        
		10'h176:out <=8'b00001100;        
		10'h177:out <=8'b00000000;        
		10'h178:out <=8'b00000000;        // /
		10'h179:out <=8'b00000001;        
		10'h17A:out <=8'b00000010;        
		10'h17B:out <=8'b00000100;        
		10'h17C:out <=8'b00001000;        
		10'h17D:out <=8'b00010000;        
		10'h17E:out <=8'b00000000;        
		10'h17F:out <=8'b00000000;        
		10'h180:out <=8'b00001110;        // 0
		10'h181:out <=8'b00010001;        
		10'h182:out <=8'b00010011;        
		10'h183:out <=8'b00010101;        
		10'h184:out <=8'b00011001;        
		10'h185:out <=8'b00010001;        
		10'h186:out <=8'b00001110;        
		10'h187:out <=8'b00000000;        
		10'h188:out <=8'b00000100;        // 1
		10'h189:out <=8'b00001100;        
		10'h18A:out <=8'b00000100;        
		10'h18B:out <=8'b00000100;        
		10'h18C:out <=8'b00000100;        
		10'h18D:out <=8'b00000100;        
		10'h18E:out <=8'b00001110;        
		10'h18F:out <=8'b00000000;        
		10'h190:out <=8'b00001110;        // 2
		10'h191:out <=8'b00010001;        
		10'h192:out <=8'b00000001;        
		10'h193:out <=8'b00000010;        
		10'h194:out <=8'b00000100;        
		10'h195:out <=8'b00001000;        
		10'h196:out <=8'b00011111;        
		10'h197:out <=8'b00000000;        
		10'h198:out <=8'b00011111;        // 3
		10'h199:out <=8'b00000010;        
		10'h19A:out <=8'b00000100;        
		10'h19B:out <=8'b00000010;        
		10'h19C:out <=8'b00000001;        
		10'h19D:out <=8'b00010001;        
		10'h19E:out <=8'b00001110;        
		10'h19F:out <=8'b00000000;        
		10'h1A0:out <=8'b00000010;        // 4
		10'h1A1:out <=8'b00000110;        
		10'h1A2:out <=8'b00001010;        
		10'h1A3:out <=8'b00010010;        
		10'h1A4:out <=8'b00011111;        
		10'h1A5:out <=8'b00000010;        
		10'h1A6:out <=8'b00000010;        
		10'h1A7:out <=8'b00000000;        
		10'h1A8:out <=8'b00011111;        // 5
		10'h1A9:out <=8'b00010000;        
		10'h1AA:out <=8'b00011110;        
		10'h1AB:out <=8'b00000001;        
		10'h1AC:out <=8'b00000001;        
		10'h1AD:out <=8'b00010001;        
		10'h1AE:out <=8'b00001110;        
		10'h1AF:out <=8'b00000000;        
		10'h1B0:out <=8'b00000110;        // 6
		10'h1B1:out <=8'b00001000;        
		10'h1B2:out <=8'b00010000;        
		10'h1B3:out <=8'b00011110;        
		10'h1B4:out <=8'b00010001;        
		10'h1B5:out <=8'b00010001;        
		10'h1B6:out <=8'b00001110;        
		10'h1B7:out <=8'b00000000;        
		10'h1B8:out <=8'b00011111;        // 7
		10'h1B9:out <=8'b00000001;        
		10'h1BA:out <=8'b00000010;        
		10'h1BB:out <=8'b00000100;        
		10'h1BC:out <=8'b00000100;        
		10'h1BD:out <=8'b00000100;        
		10'h1BE:out <=8'b00000100;        
		10'h1BF:out <=8'b00000000;        
		10'h1C0:out <=8'b00011110;        // 8
		10'h1C1:out <=8'b00010001;        
		10'h1C2:out <=8'b00010001;        
		10'h1C3:out <=8'b00001110;        
		10'h1C4:out <=8'b00010001;        
		10'h1C5:out <=8'b00010001;        
		10'h1C6:out <=8'b00001110;        
		10'h1C7:out <=8'b00000000;        
		10'h1C8:out <=8'b00001110;        // 9
		10'h1C9:out <=8'b00010001;        
		10'h1CA:out <=8'b00010001;        
		10'h1CB:out <=8'b00001111;        
		10'h1CC:out <=8'b00000001;        
		10'h1CD:out <=8'b00000010;        
		10'h1CE:out <=8'b00001100;        
		10'h1CF:out <=8'b00000000;        
		10'h1D0:out <=8'b00000000;        // :
		10'h1D1:out <=8'b00001100;        
		10'h1D2:out <=8'b00001100;        
		10'h1D3:out <=8'b00000000;        
		10'h1D4:out <=8'b00001100;        
		10'h1D5:out <=8'b00001100;        
		10'h1D6:out <=8'b00000000;        
		10'h1D7:out <=8'b00000000;        
		10'h1D8:out <=8'b00000000;        // ;
		10'h1D9:out <=8'b00001100;        
		10'h1DA:out <=8'b00001100;        
		10'h1DB:out <=8'b00000000;        
		10'h1DC:out <=8'b00001100;        
		10'h1DD:out <=8'b00000100;        
		10'h1DE:out <=8'b00001000;        
		10'h1DF:out <=8'b00000000;        
		10'h1E0:out <=8'b00000010;        // <
		10'h1E1:out <=8'b00000100;        
		10'h1E2:out <=8'b00001000;        
		10'h1E3:out <=8'b00010000;        
		10'h1E4:out <=8'b00001000;        
		10'h1E5:out <=8'b00000100;        
		10'h1E6:out <=8'b00000010;        
		10'h1E7:out <=8'b00000000;        
		10'h1E8:out <=8'b00000000;        // =
		10'h1E9:out <=8'b00000000;        
		10'h1EA:out <=8'b00011111;        
		10'h1EB:out <=8'b00000000;        
		10'h1EC:out <=8'b00011111;        
		10'h1ED:out <=8'b00000000;        
		10'h1EE:out <=8'b00000000;        
		10'h1EF:out <=8'b00000000;        
		10'h1F0:out <=8'b00001000;        // >
		10'h1F1:out <=8'b00000100;        
		10'h1F2:out <=8'b00000010;        
		10'h1F3:out <=8'b00000001;        
		10'h1F4:out <=8'b00000010;        
		10'h1F5:out <=8'b00000100;        
		10'h1F6:out <=8'b00001000;        
		10'h1F7:out <=8'b00000000;        
		10'h1F8:out <=8'b00001110;        // ?
		10'h1F9:out <=8'b00010001;        
		10'h1FA:out <=8'b00000001;        
		10'h1FB:out <=8'b00000010;        
		10'h1FC:out <=8'b00000100;        
		10'h1FD:out <=8'b00000000;        
		10'h1FE:out <=8'b00000100;        
		10'h1FF:out <=8'b00000000;        
		10'h200:out <=8'b00001110;        // @
		10'h201:out <=8'b00010001;        
		10'h202:out <=8'b00000001;        
		10'h203:out <=8'b00001101;        
		10'h204:out <=8'b00010101;        
		10'h205:out <=8'b00010101;        
		10'h206:out <=8'b00001110;        
		10'h207:out <=8'b00000000;        
		10'h208:out <=8'b00001110;        // A
		10'h209:out <=8'b00010001;        
		10'h20A:out <=8'b00010001;        
		10'h20B:out <=8'b00010001;        
		10'h20C:out <=8'b00011111;        
		10'h20D:out <=8'b00010001;        
		10'h20E:out <=8'b00010001;        
		10'h20F:out <=8'b00000000;        
		10'h210:out <=8'b00011110;        // B
		10'h211:out <=8'b00001001;        
		10'h212:out <=8'b00001001;        
		10'h213:out <=8'b00001110;        
		10'h214:out <=8'b00001001;        
		10'h215:out <=8'b00001001;        
		10'h216:out <=8'b00011110;        
		10'h217:out <=8'b00000000;        
		10'h218:out <=8'b00001110;        // C
		10'h219:out <=8'b00010001;        
		10'h21A:out <=8'b00010000;        
		10'h21B:out <=8'b00010000;        
		10'h21C:out <=8'b00010000;        
		10'h21D:out <=8'b00010001;        
		10'h21E:out <=8'b00001110;        
		10'h21F:out <=8'b00000000;        
		10'h220:out <=8'b00011110;        // D
		10'h221:out <=8'b00001001;        
		10'h222:out <=8'b00001001;        
		10'h223:out <=8'b00001001;        
		10'h224:out <=8'b00001001;        
		10'h225:out <=8'b00001001;        
		10'h226:out <=8'b00011110;        
		10'h227:out <=8'b00000000;        
		10'h228:out <=8'b00011111;        // E
		10'h229:out <=8'b00010000;        
		10'h22A:out <=8'b00010000;        
		10'h22B:out <=8'b00011111;        
		10'h22C:out <=8'b00010000;        
		10'h22D:out <=8'b00010000;        
		10'h22E:out <=8'b00011111;        
		10'h22F:out <=8'b00000000;        
		10'h230:out <=8'b00011111;        // F
		10'h231:out <=8'b00010000;        
		10'h232:out <=8'b00010000;        
		10'h233:out <=8'b00011110;        
		10'h234:out <=8'b00010000;        
		10'h235:out <=8'b00010000;        
		10'h236:out <=8'b00010000;        
		10'h237:out <=8'b00000000;        
		10'h238:out <=8'b00001110;        // G
		10'h239:out <=8'b00010001;        
		10'h23A:out <=8'b00010000;        
		10'h23B:out <=8'b00010011;        
		10'h23C:out <=8'b00010001;        
		10'h23D:out <=8'b00010001;        
		10'h23E:out <=8'b00001111;        
		10'h23F:out <=8'b00000000;        
		10'h240:out <=8'b00010001;        // H
		10'h241:out <=8'b00010001;        
		10'h242:out <=8'b00010001;        
		10'h243:out <=8'b00011111;        
		10'h244:out <=8'b00010001;        
		10'h245:out <=8'b00010001;        
		10'h246:out <=8'b00010001;        
		10'h247:out <=8'b00000000;        
		10'h248:out <=8'b00001110;        // I
		10'h249:out <=8'b00000100;        
		10'h24A:out <=8'b00000100;        
		10'h24B:out <=8'b00000100;        
		10'h24C:out <=8'b00000100;        
		10'h24D:out <=8'b00000100;        
		10'h24E:out <=8'b00001110;        
		10'h24F:out <=8'b00000000;        
		10'h250:out <=8'b00000111;        // J
		10'h251:out <=8'b00000010;        
		10'h252:out <=8'b00000010;        
		10'h253:out <=8'b00000010;        
		10'h254:out <=8'b00000010;        
		10'h255:out <=8'b00010010;        
		10'h256:out <=8'b00001100;        
		10'h257:out <=8'b00000000;        
		10'h258:out <=8'b00010001;        // K
		10'h259:out <=8'b00010010;        
		10'h25A:out <=8'b00010100;        
		10'h25B:out <=8'b00011000;        
		10'h25C:out <=8'b00010100;        
		10'h25D:out <=8'b00010010;        
		10'h25E:out <=8'b00010001;        
		10'h25F:out <=8'b00000000;        
		10'h260:out <=8'b00010000;        // L
		10'h261:out <=8'b00010000;        
		10'h262:out <=8'b00010000;        
		10'h263:out <=8'b00010000;        
		10'h264:out <=8'b00010000;        
		10'h265:out <=8'b00010000;        
		10'h266:out <=8'b00011111;        
		10'h267:out <=8'b00000000;        
		10'h268:out <=8'b00010001;        // M
		10'h269:out <=8'b00011011;        
		10'h26A:out <=8'b00010101;        
		10'h26B:out <=8'b00010101;        
		10'h26C:out <=8'b00010001;        
		10'h26D:out <=8'b00010001;        
		10'h26E:out <=8'b00010001;        
		10'h26F:out <=8'b00000000;        
		10'h270:out <=8'b00010001;        // N
		10'h271:out <=8'b00011001;        
		10'h272:out <=8'b00011001;        
		10'h273:out <=8'b00010101;        
		10'h274:out <=8'b00010011;        
		10'h275:out <=8'b00010011;        
		10'h276:out <=8'b00010001;        
		10'h277:out <=8'b00000000;        
		10'h278:out <=8'b00001110;        // O
		10'h279:out <=8'b00010001;        
		10'h27A:out <=8'b00010001;        
		10'h27B:out <=8'b00010001;        
		10'h27C:out <=8'b00010001;        
		10'h27D:out <=8'b00010001;        
		10'h27E:out <=8'b00001110;        
		10'h27F:out <=8'b00000000;        
		10'h280:out <=8'b00011110;        // P
		10'h281:out <=8'b00010001;        
		10'h282:out <=8'b00010001;        
		10'h283:out <=8'b00011110;        
		10'h284:out <=8'b00010000;        
		10'h285:out <=8'b00010000;        
		10'h286:out <=8'b00010000;        
		10'h287:out <=8'b00000000;        
		10'h288:out <=8'b00001110;        // Q
		10'h289:out <=8'b00010001;        
		10'h28A:out <=8'b00010001;        
		10'h28B:out <=8'b00010001;        
		10'h28C:out <=8'b00010101;        
		10'h28D:out <=8'b00010010;        
		10'h28E:out <=8'b00011101;        
		10'h28F:out <=8'b00000000;        
		10'h290:out <=8'b00011110;        // R
		10'h291:out <=8'b00010001;        
		10'h292:out <=8'b00010001;        
		10'h293:out <=8'b00011110;        
		10'h294:out <=8'b00010100;        
		10'h295:out <=8'b00010010;        
		10'h296:out <=8'b00010001;        
		10'h297:out <=8'b00000000;        
		10'h298:out <=8'b00001110;        // S
		10'h299:out <=8'b00010001;        
		10'h29A:out <=8'b00010000;        
		10'h29B:out <=8'b00001110;        
		10'h29C:out <=8'b00000001;        
		10'h29D:out <=8'b00010001;        
		10'h29E:out <=8'b00001110;        
		10'h29F:out <=8'b00000000;        
		10'h2A0:out <=8'b00011111;        // T
		10'h2A1:out <=8'b00000100;        
		10'h2A2:out <=8'b00000100;        
		10'h2A3:out <=8'b00000100;        
		10'h2A4:out <=8'b00000100;        
		10'h2A5:out <=8'b00000100;        
		10'h2A6:out <=8'b00000100;        
		10'h2A7:out <=8'b00000000;        
		10'h2A8:out <=8'b00010001;        // U
		10'h2A9:out <=8'b00010001;        
		10'h2AA:out <=8'b00010001;        
		10'h2AB:out <=8'b00010001;        
		10'h2AC:out <=8'b00010001;        
		10'h2AD:out <=8'b00010001;        
		10'h2AE:out <=8'b00001110;        
		10'h2AF:out <=8'b00000000;        
		10'h2B0:out <=8'b00010001;        // V
		10'h2B1:out <=8'b00010001;        
		10'h2B2:out <=8'b00010001;        
		10'h2B3:out <=8'b00010001;        
		10'h2B4:out <=8'b00010001;        
		10'h2B5:out <=8'b00001010;        
		10'h2B6:out <=8'b00000100;        
		10'h2B7:out <=8'b00000000;        
		10'h2B8:out <=8'b00010001;        // W
		10'h2B9:out <=8'b00010001;        
		10'h2BA:out <=8'b00010001;        
		10'h2BB:out <=8'b00010101;        
		10'h2BC:out <=8'b00010101;        
		10'h2BD:out <=8'b00011011;        
		10'h2BE:out <=8'b00010001;        
		10'h2BF:out <=8'b00000000;        
		10'h2C0:out <=8'b00010001;        // X
		10'h2C1:out <=8'b00010001;        
		10'h2C2:out <=8'b00001010;        
		10'h2C3:out <=8'b00000100;        
		10'h2C4:out <=8'b00001010;        
		10'h2C5:out <=8'b00010001;        
		10'h2C6:out <=8'b00010001;        
		10'h2C7:out <=8'b00000000;        
		10'h2C8:out <=8'b00010001;        // Y
		10'h2C9:out <=8'b00010001;        
		10'h2CA:out <=8'b00010001;        
		10'h2CB:out <=8'b00001010;        
		10'h2CC:out <=8'b00000100;        
		10'h2CD:out <=8'b00000100;        
		10'h2CE:out <=8'b00000100;        
		10'h2CF:out <=8'b00000000;        
		10'h2D0:out <=8'b00011111;        // Z
		10'h2D1:out <=8'b00000001;        
		10'h2D2:out <=8'b00000010;        
		10'h2D3:out <=8'b00000100;        
		10'h2D4:out <=8'b00001000;        
		10'h2D5:out <=8'b00010000;        
		10'h2D6:out <=8'b00011111;        
		10'h2D7:out <=8'b00000000;        
		10'h2D8:out <=8'b00001110;        // [
		10'h2D9:out <=8'b00001000;        
		10'h2DA:out <=8'b00001000;        
		10'h2DB:out <=8'b00001000;        
		10'h2DC:out <=8'b00001000;        
		10'h2DD:out <=8'b00001000;        
		10'h2DE:out <=8'b00001110;        
		10'h2DF:out <=8'b00000000;        
		10'h2E0:out <=8'b00000000;        // \
		10'h2E1:out <=8'b00010000;        
		10'h2E2:out <=8'b00001000;        
		10'h2E3:out <=8'b00000100;        
		10'h2E4:out <=8'b00000010;        
		10'h2E5:out <=8'b00000001;        
		10'h2E6:out <=8'b00000000;        
		10'h2E7:out <=8'b00000000;        
		10'h2E8:out <=8'b00001110;        // ]
		10'h2E9:out <=8'b00000010;        
		10'h2EA:out <=8'b00000010;        
		10'h2EB:out <=8'b00000010;        
		10'h2EC:out <=8'b00000010;        
		10'h2ED:out <=8'b00000010;        
		10'h2EE:out <=8'b00001110;        
		10'h2EF:out <=8'b00000000;        
		10'h2F0:out <=8'b00000100;        // ^
		10'h2F1:out <=8'b00001010;        
		10'h2F2:out <=8'b00010001;        
		10'h2F3:out <=8'b00000000;        
		10'h2F4:out <=8'b00000000;        
		10'h2F5:out <=8'b00000000;        
		10'h2F6:out <=8'b00000000;        
		10'h2F7:out <=8'b00000000;        
		10'h2F8:out <=8'b00000000;        // _
		10'h2F9:out <=8'b00000000;        
		10'h2FA:out <=8'b00000000;        
		10'h2FB:out <=8'b00000000;        
		10'h2FC:out <=8'b00000000;        
		10'h2FD:out <=8'b00000000;        
		10'h2FE:out <=8'b00011111;        
		10'h2FF:out <=8'b00000000;        
		10'h300:out <=8'b00010000;        // `
		10'h301:out <=8'b00001000;        
		10'h302:out <=8'b00000100;        
		10'h303:out <=8'b00000000;        
		10'h304:out <=8'b00000000;        
		10'h305:out <=8'b00000000;        
		10'h306:out <=8'b00000000;        
		10'h307:out <=8'b00000000;        
		10'h308:out <=8'b00000000;        // a
		10'h309:out <=8'b00000000;        
		10'h30A:out <=8'b00001110;        
		10'h30B:out <=8'b00000001;        
		10'h30C:out <=8'b00001111;        
		10'h30D:out <=8'b00010001;        
		10'h30E:out <=8'b00001111;        
		10'h30F:out <=8'b00000000;        
		10'h310:out <=8'b00010000;        // b
		10'h311:out <=8'b00010000;        
		10'h312:out <=8'b00010110;        
		10'h313:out <=8'b00011001;        
		10'h314:out <=8'b00010001;        
		10'h315:out <=8'b00010001;        
		10'h316:out <=8'b00011110;        
		10'h317:out <=8'b00000000;        
		10'h318:out <=8'b00000000;        // c
		10'h319:out <=8'b00000000;        
		10'h31A:out <=8'b00001110;        
		10'h31B:out <=8'b00010001;        
		10'h31C:out <=8'b00010000;        
		10'h31D:out <=8'b00010001;        
		10'h31E:out <=8'b00001110;        
		10'h31F:out <=8'b00000000;        
		10'h320:out <=8'b00000001;        // d
		10'h321:out <=8'b00000001;        
		10'h322:out <=8'b00001101;        
		10'h323:out <=8'b00010011;        
		10'h324:out <=8'b00010001;        
		10'h325:out <=8'b00010001;        
		10'h326:out <=8'b00001111;        
		10'h327:out <=8'b00000000;        
		10'h328:out <=8'b00000000;        // e
		10'h329:out <=8'b00000000;        
		10'h32A:out <=8'b00001110;        
		10'h32B:out <=8'b00010001;        
		10'h32C:out <=8'b00011111;        
		10'h32D:out <=8'b00010000;        
		10'h32E:out <=8'b00001110;        
		10'h32F:out <=8'b00000000;        
		10'h330:out <=8'b00000010;        // f
		10'h331:out <=8'b00000101;        
		10'h332:out <=8'b00000100;        
		10'h333:out <=8'b00001110;        
		10'h334:out <=8'b00000100;        
		10'h335:out <=8'b00000100;        
		10'h336:out <=8'b00000100;        
		10'h337:out <=8'b00000000;        
		10'h338:out <=8'b00000000;        // g
		10'h339:out <=8'b00001101;        
		10'h33A:out <=8'b00010011;        
		10'h33B:out <=8'b00010011;        
		10'h33C:out <=8'b00001101;        
		10'h33D:out <=8'b00000001;        
		10'h33E:out <=8'b00001110;        
		10'h33F:out <=8'b00000000;        
		10'h340:out <=8'b00010000;        // h
		10'h341:out <=8'b00010000;        
		10'h342:out <=8'b00010110;        
		10'h343:out <=8'b00011001;        
		10'h344:out <=8'b00010001;        
		10'h345:out <=8'b00010001;        
		10'h346:out <=8'b00010001;        
		10'h347:out <=8'b00000000;        
		10'h348:out <=8'b00000100;        // i
		10'h349:out <=8'b00000000;        
		10'h34A:out <=8'b00001100;        
		10'h34B:out <=8'b00000100;        
		10'h34C:out <=8'b00000100;        
		10'h34D:out <=8'b00000100;        
		10'h34E:out <=8'b00001110;        
		10'h34F:out <=8'b00000000;        
		10'h350:out <=8'b00000010;        // j
		10'h351:out <=8'b00000000;        
		10'h352:out <=8'b00000110;        
		10'h353:out <=8'b00000010;        
		10'h354:out <=8'b00000010;        
		10'h355:out <=8'b00010010;        
		10'h356:out <=8'b00001100;        
		10'h357:out <=8'b00000000;        
		10'h358:out <=8'b00001000;        // k
		10'h359:out <=8'b00001000;        
		10'h35A:out <=8'b00001001;        
		10'h35B:out <=8'b00001010;        
		10'h35C:out <=8'b00001100;        
		10'h35D:out <=8'b00001010;        
		10'h35E:out <=8'b00001001;        
		10'h35F:out <=8'b00000000;        
		10'h360:out <=8'b00001100;        // l
		10'h361:out <=8'b00000100;        
		10'h362:out <=8'b00000100;        
		10'h363:out <=8'b00000100;        
		10'h364:out <=8'b00000100;        
		10'h365:out <=8'b00000100;        
		10'h366:out <=8'b00001110;        
		10'h367:out <=8'b00000000;        
		10'h368:out <=8'b00000000;        // m
		10'h369:out <=8'b00000000;        
		10'h36A:out <=8'b00011010;        
		10'h36B:out <=8'b00010101;        
		10'h36C:out <=8'b00010101;        
		10'h36D:out <=8'b00010101;        
		10'h36E:out <=8'b00010101;        
		10'h36F:out <=8'b00000000;        
		10'h370:out <=8'b00000000;        // n
		10'h371:out <=8'b00000000;        
		10'h372:out <=8'b00010110;        
		10'h373:out <=8'b00011001;        
		10'h374:out <=8'b00010001;        
		10'h375:out <=8'b00010001;        
		10'h376:out <=8'b00010001;        
		10'h377:out <=8'b00000000;        
		10'h378:out <=8'b00000000;        // o
		10'h379:out <=8'b00000000;        
		10'h37A:out <=8'b00001110;        
		10'h37B:out <=8'b00010001;        
		10'h37C:out <=8'b00010001;        
		10'h37D:out <=8'b00010001;        
		10'h37E:out <=8'b00001110;        
		10'h37F:out <=8'b00000000;        
		10'h380:out <=8'b00000000;        // p
		10'h381:out <=8'b00010110;        
		10'h382:out <=8'b00011001;        
		10'h383:out <=8'b00011001;        
		10'h384:out <=8'b00010110;        
		10'h385:out <=8'b00010000;        
		10'h386:out <=8'b00010000;        
		10'h387:out <=8'b00000000;        
		10'h388:out <=8'b00000000;        // q
		10'h389:out <=8'b00001101;        
		10'h38A:out <=8'b00010011;        
		10'h38B:out <=8'b00010011;        
		10'h38C:out <=8'b00001101;        
		10'h38D:out <=8'b00000001;        
		10'h38E:out <=8'b00000001;        
		10'h38F:out <=8'b00000000;        
		10'h390:out <=8'b00000000;        // r
		10'h391:out <=8'b00000000;        
		10'h392:out <=8'b00010110;        
		10'h393:out <=8'b00011001;        
		10'h394:out <=8'b00010000;        
		10'h395:out <=8'b00010000;        
		10'h396:out <=8'b00010000;        
		10'h397:out <=8'b00000000;        
		10'h398:out <=8'b00000000;        // s
		10'h399:out <=8'b00000000;        
		10'h39A:out <=8'b00001111;        
		10'h39B:out <=8'b00010000;        
		10'h39C:out <=8'b00011110;        
		10'h39D:out <=8'b00000001;        
		10'h39E:out <=8'b00011111;        
		10'h39F:out <=8'b00000000;        
		10'h3A0:out <=8'b00001000;        // t
		10'h3A1:out <=8'b00001000;        
		10'h3A2:out <=8'b00011100;        
		10'h3A3:out <=8'b00001000;        
		10'h3A4:out <=8'b00001000;        
		10'h3A5:out <=8'b00001001;        
		10'h3A6:out <=8'b00000110;        
		10'h3A7:out <=8'b00000000;        
		10'h3A8:out <=8'b00000000;        // u
		10'h3A9:out <=8'b00000000;        
		10'h3AA:out <=8'b00010010;        
		10'h3AB:out <=8'b00010010;        
		10'h3AC:out <=8'b00010010;        
		10'h3AD:out <=8'b00010010;        
		10'h3AE:out <=8'b00001101;        
		10'h3AF:out <=8'b00000000;        
		10'h3B0:out <=8'b00000000;        // v
		10'h3B1:out <=8'b00000000;        
		10'h3B2:out <=8'b00010001;        
		10'h3B3:out <=8'b00010001;        
		10'h3B4:out <=8'b00010001;        
		10'h3B5:out <=8'b00001010;        
		10'h3B6:out <=8'b00000100;        
		10'h3B7:out <=8'b00000000;        
		10'h3B8:out <=8'b00000000;        // w
		10'h3B9:out <=8'b00000000;        
		10'h3BA:out <=8'b00010001;        
		10'h3BB:out <=8'b00010001;        
		10'h3BC:out <=8'b00010101;        
		10'h3BD:out <=8'b00010101;        
		10'h3BE:out <=8'b00001010;        
		10'h3BF:out <=8'b00000000;        
		10'h3C0:out <=8'b00000000;        // x
		10'h3C1:out <=8'b00000000;        
		10'h3C2:out <=8'b00010001;        
		10'h3C3:out <=8'b00001010;        
		10'h3C4:out <=8'b00000100;        
		10'h3C5:out <=8'b00001010;        
		10'h3C6:out <=8'b00010001;        
		10'h3C7:out <=8'b00000000;        
		10'h3C8:out <=8'b00000000;        // y
		10'h3C9:out <=8'b00000000;        
		10'h3CA:out <=8'b00010001;        
		10'h3CB:out <=8'b00010001;        
		10'h3CC:out <=8'b00010011;        
		10'h3CD:out <=8'b00001101;        
		10'h3CE:out <=8'b00000001;        
		10'h3CF:out <=8'b00001110;        
		10'h3D0:out <=8'b00000000;        // z
		10'h3D1:out <=8'b00000000;        
		10'h3D2:out <=8'b00011111;        
		10'h3D3:out <=8'b00000010;        
		10'h3D4:out <=8'b00000100;        
		10'h3D5:out <=8'b00001000;        
		10'h3D6:out <=8'b00011111;        
		10'h3D7:out <=8'b00000000;        
		10'h3D8:out <=8'b00000010;        // {
		10'h3D9:out <=8'b00000100;        
		10'h3DA:out <=8'b00000100;        
		10'h3DB:out <=8'b00001000;        
		10'h3DC:out <=8'b00000100;        
		10'h3DD:out <=8'b00000100;        
		10'h3DE:out <=8'b00000010;        
		10'h3DF:out <=8'b00000000;        
		10'h3E0:out <=8'b00000100;        // |
		10'h3E1:out <=8'b00000100;        
		10'h3E2:out <=8'b00000100;        
		10'h3E3:out <=8'b00000000;        
		10'h3E4:out <=8'b00000100;        
		10'h3E5:out <=8'b00000100;        
		10'h3E6:out <=8'b00000100;        
		10'h3E7:out <=8'b00000000;        
		10'h3E8:out <=8'b00001000;        // }
		10'h3E9:out <=8'b00000100;        
		10'h3EA:out <=8'b00000100;        
		10'h3EB:out <=8'b00000010;        
		10'h3EC:out <=8'b00000100;        
		10'h3ED:out <=8'b00000100;        
		10'h3EE:out <=8'b00001000;        
		10'h3EF:out <=8'b00000000;        
		10'h3F0:out <=8'b00001000;        // ~
		10'h3F1:out <=8'b00010101;        
		10'h3F2:out <=8'b00000010;        
		10'h3F3:out <=8'b00000000;        
		10'h3F4:out <=8'b00000000;        
		10'h3F5:out <=8'b00000000;        
		10'h3F6:out <=8'b00000000;        
		10'h3F7:out <=8'b00000000;               
    default : out <= 0;
  endcase
end
endmodule

//DEC 	OCT 	HEX 	BIN 	Symbol 	HTML Number 	HTML Name 	Description
//0	000	00	00000000	NUL	&#000;	 	Null char
//1	001	01	00000001	SOH	&#001;	 	Start of Heading
//2	002	02	00000010	STX	&#002;	 	Start of Text
//3	003	03	00000011	ETX	&#003;	 	End of Text
//4	004	04	00000100	EOT	&#004;	 	End of Transmission
//5	005	05	00000101	ENQ	&#005;	 	Enquiry
//6	006	06	00000110	ACK	&#006;	 	Acknowledgment
//7	007	07	00000111	BEL	&#007;	 	Bell
//8	010	08	00001000	BS	&#008;	 	Back Space
//9	011	09	00001001	HT	&#009;	 	Horizontal Tab
//10	012	0A	00001010	LF	&#010;	 	Line Feed
//11	013	0B	00001011	VT	&#011;	 	Vertical Tab
//12	014	0C	00001100	FF	&#012;	 	Form Feed
//13	015	0D	00001101	CR	&#013;	 	Carriage Return
//14	016	0E	00001110	SO	&#014;	 	Shift Out / X-On
//15	017	0F	00001111	SI	&#015;	 	Shift In / X-Off
//16	020	10	00010000	DLE	&#016;	 	Data Line Escape
//17	021	11	00010001	DC1	&#017;	 	Device Control 1 (oft. XON)
//18	022	12	00010010	DC2	&#018;	 	Device Control 2
//19	023	13	00010011	DC3	&#019;	 	Device Control 3 (oft. XOFF)
//20	024	14	00010100	DC4	&#020;	 	Device Control 4
//21	025	15	00010101	NAK	&#021;	 	Negative Acknowledgement
//22	026	16	00010110	SYN	&#022;	 	Synchronous Idle
//23	027	17	00010111	ETB	&#023;	 	End of Transmit Block
//24	030	18	00011000	CAN	&#024;	 	Cancel
//25	031	19	00011001	EM	&#025;	 	End of Medium
//26	032	1A	00011010	SUB	&#026;	 	Substitute
//27	033	1B	00011011	ESC	&#027;	 	Escape
//28	034	1C	00011100	FS	&#028;	 	File Separator
//29	035	1D	00011101	GS	&#029;	 	Group Separator
//30	036	1E	00011110	RS	&#030;	 	Record Separator
//31	037	1F	00011111	US	&#031;	 	Unit Separator
//32	040	20	00100000	 	&#32;	 	Space
//33	041	21	00100001	!	&#33;	 	Exclamation mark
//34	042	22	00100010	"	&#34;	&quot;	Double quotes (or speech marks)
//35	043	23	00100011	#	&#35;	 	Number
//36	044	24	00100100	$	&#36;	 	Dollar
//37	045	25	00100101	%	&#37;	 	Procenttecken
//38	046	26	00100110	&	&#38;	&amp;	Ampersand
//39	047	27	00100111	'	&#39;	 	Single quote
//40	050	28	00101000	(	&#40;	 	Open parenthesis (or open bracket)
//41	051	29	00101001	)	&#41;	 	Close parenthesis (or close bracket)
//42	052	2A	00101010	*	&#42;	 	Asterisk
//43	053	2B	00101011	+	&#43;	 	Plus
//44	054	2C	00101100	,	&#44;	 	Comma
//45	055	2D	00101101	-	&#45;	 	Hyphen
//46	056	2E	00101110	.	&#46;	 	Period, dot or full stop
//47	057	2F	00101111	/	&#47;	 	Slash or divide
//48	060	30	00110000	0	&#48;	 	Zero
//49	061	31	00110001	1	&#49;	 	One
//50	062	32	00110010	2	&#50;	 	Two
//51	063	33	00110011	3	&#51;	 	Three
//52	064	34	00110100	4	&#52;	 	Four
//53	065	35	00110101	5	&#53;	 	Five
//54	066	36	00110110	6	&#54;	 	Six
//55	067	37	00110111	7	&#55;	 	Seven
//56	070	38	00111000	8	&#56;	 	Eight
//57	071	39	00111001	9	&#57;	 	Nine
//58	072	3A	00111010	:	&#58;	 	Colon
//59	073	3B	00111011	;	&#59;	 	Semicolon
//60	074	3C	00111100	<	&#60;	&lt;	Less than (or open angled bracket)
//61	075	3D	00111101	=	&#61;	 	Equals
//62	076	3E	00111110	>	&#62;	&gt;	Greater than (or close angled bracket)
//63	077	3F	00111111	?	&#63;	 	Question mark
//64	100	40	01000000	@	&#64;	 	At symbol
//65	101	41	01000001	A	&#65;	 	Uppercase A
//66	102	42	01000010	B	&#66;	 	Uppercase B
//67	103	43	01000011	C	&#67;	 	Uppercase C
//68	104	44	01000100	D	&#68;	 	Uppercase D
//69	105	45	01000101	E	&#69;	 	Uppercase E
//70	106	46	01000110	F	&#70;	 	Uppercase F
//71	107	47	01000111	G	&#71;	 	Uppercase G
//72	110	48	01001000	H	&#72;	 	Uppercase H
//73	111	49	01001001	I	&#73;	 	Uppercase I
//74	112	4A	01001010	J	&#74;	 	Uppercase J
//75	113	4B	01001011	K	&#75;	 	Uppercase K
//76	114	4C	01001100	L	&#76;	 	Uppercase L
//77	115	4D	01001101	M	&#77;	 	Uppercase M
//78	116	4E	01001110	N	&#78;	 	Uppercase N
//79	117	4F	01001111	O	&#79;	 	Uppercase O
//80	120	50	01010000	P	&#80;	 	Uppercase P
//81	121	51	01010001	Q	&#81;	 	Uppercase Q
//82	122	52	01010010	R	&#82;	 	Uppercase R
//83	123	53	01010011	S	&#83;	 	Uppercase S
//84	124	54	01010100	T	&#84;	 	Uppercase T
//85	125	55	01010101	U	&#85;	 	Uppercase U
//86	126	56	01010110	V	&#86;	 	Uppercase V
//87	127	57	01010111	W	&#87;	 	Uppercase W
//88	130	58	01011000	X	&#88;	 	Uppercase X
//89	131	59	01011001	Y	&#89;	 	Uppercase Y
//90	132	5A	01011010	Z	&#90;	 	Uppercase Z
//91	133	5B	01011011	[	&#91;	 	Opening bracket
//92	134	5C	01011100	\	&#92;	 	Backslash
//93	135	5D	01011101	]	&#93;	 	Closing bracket
//94	136	5E	01011110	^	&#94;	 	Caret - circumflex
//95	137	5F	01011111	_	&#95;	 	Underscore
//96	140	60	01100000	`	&#96;	 	Grave accent
//97	141	61	01100001	a	&#97;	 	Lowercase a
//98	142	62	01100010	b	&#98;	 	Lowercase b
//99	143	63	01100011	c	&#99;	 	Lowercase c
//100	144	64	01100100	d	&#100;	 	Lowercase d
//101	145	65	01100101	e	&#101;	 	Lowercase e
//102	146	66	01100110	f	&#102;	 	Lowercase f
//103	147	67	01100111	g	&#103;	 	Lowercase g
//104	150	68	01101000	h	&#104;	 	Lowercase h
//105	151	69	01101001	i	&#105;	 	Lowercase i
//106	152	6A	01101010	j	&#106;	 	Lowercase j
//107	153	6B	01101011	k	&#107;	 	Lowercase k
//108	154	6C	01101100	l	&#108;	 	Lowercase l
//109	155	6D	01101101	m	&#109;	 	Lowercase m
//110	156	6E	01101110	n	&#110;	 	Lowercase n
//111	157	6F	01101111	o	&#111;	 	Lowercase o
//112	160	70	01110000	p	&#112;	 	Lowercase p
//113	161	71	01110001	q	&#113;	 	Lowercase q
//114	162	72	01110010	r	&#114;	 	Lowercase r
//115	163	73	01110011	s	&#115;	 	Lowercase s
//116	164	74	01110100	t	&#116;	 	Lowercase t
//117	165	75	01110101	u	&#117;	 	Lowercase u
//118	166	76	01110110	v	&#118;	 	Lowercase v
//119	167	77	01110111	w	&#119;	 	Lowercase w
//120	170	78	01111000	x	&#120;	 	Lowercase x
//121	171	79	01111001	y	&#121;	 	Lowercase y
//122	172	7A	01111010	z	&#122;	 	Lowercase z
//123	173	7B	01111011	{	&#123;	 	Opening brace
//124	174	7C	01111100	|	&#124;	 	Vertical bar
//125	175	7D	01111101	}	&#125;	 	Closing brace
//126	176	7E	01111110	~	&#126;	 	Equivalency sign - tilde
//127	177	7F	01111111		&#127;	 	Delete
//128	200	80	10000000	€	&#128;	&euro;	Euro sign
//129	201	81	10000001	 	 	 	 
//130	202	82	10000010	‚	&#130;	&sbquo;	Single low-9 quotation mark
//131	203	83	10000011	ƒ	&#131;	&fnof;	Latin small letter f with hook
//132	204	84	10000100	„	&#132;	&bdquo;	Double low-9 quotation mark
//133	205	85	10000101	…	&#133;	&hellip;	Horizontal ellipsis
//134	206	86	10000110	†	&#134;	&dagger;	Dagger
//135	207	87	10000111	‡	&#135;	&Dagger;	Double dagger
//136	210	88	10001000	ˆ	&#136;	&circ;	Modifier letter circumflex accent
//137	211	89	10001001	‰	&#137;	&permil;	Per mille sign
//138	212	8A	10001010	Š	&#138;	&Scaron;	Latin capital letter S with caron
//139	213	8B	10001011	‹	&#139;	&lsaquo;	Single left-pointing angle quotation
//140	214	8C	10001100	Œ	&#140;	&OElig;	Latin capital ligature OE
//141	215	8D	10001101	 	 	 	 
//142	216	8E	10001110	Ž	&#142;	 	Latin captial letter Z with caron
//143	217	8F	10001111	 	 	 	 
//144	220	90	10010000	 	 	 	 
//145	221	91	10010001	‘	&#145;	&lsquo;	Left single quotation mark
//146	222	92	10010010	’	&#146;	&rsquo;	Right single quotation mark
//147	223	93	10010011	“	&#147;	&ldquo;	Left double quotation mark
//148	224	94	10010100	”	&#148;	&rdquo;	Right double quotation mark
//149	225	95	10010101	•	&#149;	&bull;	Bullet
//150	226	96	10010110	–	&#150;	&ndash;	En dash
//151	227	97	10010111	—	&#151;	&mdash;	Em dash
//152	230	98	10011000	˜	&#152;	&tilde;	Small tilde
//153	231	99	10011001	™	&#153;	&trade;	Trade mark sign
//154	232	9A	10011010	š	&#154;	&scaron;	Latin small letter S with caron
//155	233	9B	10011011	›	&#155;	&rsaquo; 	Single right-pointing angle quotation mark
//156	234	9C	10011100	œ	&#156;	&oelig;	Latin small ligature oe
//157	235	9D	10011101	 	 	 	 
//158	236	9E	10011110	ž	&#158;	 	Latin small letter z with caron
//159	237	9F	10011111	Ÿ	&#159;	&Yuml;	Latin capital letter Y with diaeresis
//160	240	A0	10100000	 	&#160;	&nbsp;	Non-breaking space
//161	241	A1	10100001	¡	&#161;	&iexcl;	Inverted exclamation mark
//162	242	A2	10100010	¢	&#162;	&cent;	Cent sign
//163	243	A3	10100011	£	&#163;	&pound;	Pound sign
//164	244	A4	10100100	¤	&#164;	&curren;	Currency sign
//165	245	A5	10100101	¥	&#165;	&yen;	Yen sign
//166	246	A6	10100110	¦	&#166;	&brvbar;	Pipe, Broken vertical bar
//167	247	A7	10100111	§	&#167;	&sect;	Section sign
//168	250	A8	10101000	¨	&#168;	&uml;	Spacing diaeresis - umlaut
//169	251	A9	10101001	©	&#169;	&copy;	Copyright sign
//170	252	AA	10101010	ª	&#170;	&ordf;	Feminine ordinal indicator
//171	253	AB	10101011	«	&#171;	&laquo;	Left double angle quotes
//172	254	AC	10101100	¬	&#172;	&not;	Not sign
//173	255	AD	10101101	­	&#173;	&shy;	Soft hyphen
//174	256	AE	10101110	®	&#174;	&reg;	Registered trade mark sign
//175	257	AF	10101111	¯	&#175;	&macr;	Spacing macron - overline
//176	260	B0	10110000	°	&#176;	&deg;	Degree sign
//177	261	B1	10110001	±	&#177;	&plusmn;	Plus-or-minus sign
//178	262	B2	10110010	²	&#178;	&sup2;	Superscript two - squared
//179	263	B3	10110011	³	&#179;	&sup3;	Superscript three - cubed
//180	264	B4	10110100	´	&#180;	&acute;	Acute accent - spacing acute
//181	265	B5	10110101	µ	&#181;	&micro;	Micro sign
//182	266	B6	10110110	¶	&#182;	&para;	Pilcrow sign - paragraph sign
//183	267	B7	10110111	·	&#183;	&middot;	Middle dot - Georgian comma
//184	270	B8	10111000	¸	&#184;	&cedil;	Spacing cedilla
//185	271	B9	10111001	¹	&#185;	&sup1;	Superscript one
//186	272	BA	10111010	º	&#186;	&ordm;	Masculine ordinal indicator
//187	273	BB	10111011	»	&#187;	&raquo;	Right double angle quotes
//188	274	BC	10111100	¼	&#188;	&frac14;	Fraction one quarter
//189	275	BD	10111101	½	&#189;	&frac12;	Fraction one half
//190	276	BE	10111110	¾	&#190;	&frac34;	Fraction three quarters
//191	277	BF	10111111	¿	&#191;	&iquest;	Inverted question mark
//192	300	C0	11000000	À	&#192;	&Agrave;	Latin capital letter A with grave
//193	301	C1	11000001	Á	&#193;	&Aacute;	Latin capital letter A with acute
//194	302	C2	11000010	Â	&#194;	&Acirc;	Latin capital letter A with circumflex
//195	303	C3	11000011	Ã	&#195;	&Atilde;	Latin capital letter A with tilde
//196	304	C4	11000100	Ä	&#196;	&Auml;	Latin capital letter A with diaeresis
//197	305	C5	11000101	Å	&#197;	&Aring;	Latin capital letter A with ring above
//198	306	C6	11000110	Æ	&#198;	&AElig;	Latin capital letter AE
//199	307	C7	11000111	Ç	&#199;	&Ccedil;	Latin capital letter C with cedilla
//200	310	C8	11001000	È	&#200;	&Egrave;	Latin capital letter E with grave
//201	311	C9	11001001	É	&#201;	&Eacute;	Latin capital letter E with acute
//202	312	CA	11001010	Ê	&#202;	&Ecirc;	Latin capital letter E with circumflex
//203	313	CB	11001011	Ë	&#203;	&Euml;	Latin capital letter E with diaeresis
//204	314	CC	11001100	Ì	&#204;	&Igrave;	Latin capital letter I with grave
//205	315	CD	11001101	Í	&#205;	&Iacute;	Latin capital letter I with acute
//206	316	CE	11001110	Î	&#206;	&Icirc;	Latin capital letter I with circumflex
//207	317	CF	11001111	Ï	&#207;	&Iuml;	Latin capital letter I with diaeresis
//208	320	D0	11010000	Ð	&#208;	&ETH;	Latin capital letter ETH
//209	321	D1	11010001	Ñ	&#209;	&Ntilde;	Latin capital letter N with tilde
//210	322	D2	11010010	Ò	&#210;	&Ograve;	Latin capital letter O with grave
//211	323	D3	11010011	Ó	&#211;	&Oacute;	Latin capital letter O with acute
//212	324	D4	11010100	Ô	&#212;	&Ocirc;	Latin capital letter O with circumflex
//213	325	D5	11010101	Õ	&#213;	&Otilde;	Latin capital letter O with tilde
//214	326	D6	11010110	Ö	&#214;	&Ouml;	Latin capital letter O with diaeresis
//215	327	D7	11010111	×	&#215;	&times;	Multiplication sign
//216	330	D8	11011000	Ø	&#216;	&Oslash;	Latin capital letter O with slash
//217	331	D9	11011001	Ù	&#217;	&Ugrave;	Latin capital letter U with grave
//218	332	DA	11011010	Ú	&#218;	&Uacute;	Latin capital letter U with acute
//219	333	DB	11011011	Û	&#219;	&Ucirc;	Latin capital letter U with circumflex
//220	334	DC	11011100	Ü	&#220;	&Uuml;	Latin capital letter U with diaeresis
//221	335	DD	11011101	Ý	&#221;	&Yacute;	Latin capital letter Y with acute
//222	336	DE	11011110	Þ	&#222;	&THORN;	Latin capital letter THORN
//223	337	DF	11011111	ß	&#223;	&szlig;	Latin small letter sharp s - ess-zed
//224	340	E0	11100000	à	&#224;	&agrave;	Latin small letter a with grave
//225	341	E1	11100001	á	&#225;	&aacute;	Latin small letter a with acute
//226	342	E2	11100010	â	&#226;	&acirc;	Latin small letter a with circumflex
//227	343	E3	11100011	ã	&#227;	&atilde;	Latin small letter a with tilde
//228	344	E4	11100100	ä	&#228;	&auml;	Latin small letter a with diaeresis
//229	345	E5	11100101	å	&#229;	&aring;	Latin small letter a with ring above
//230	346	E6	11100110	æ	&#230;	&aelig;	Latin small letter ae
//231	347	E7	11100111	ç	&#231;	&ccedil;	Latin small letter c with cedilla
//232	350	E8	11101000	è	&#232;	&egrave;	Latin small letter e with grave
//233	351	E9	11101001	é	&#233;	&eacute;	Latin small letter e with acute
//234	352	EA	11101010	ê	&#234;	&ecirc;	Latin small letter e with circumflex
//235	353	EB	11101011	ë	&#235;	&euml;	Latin small letter e with diaeresis
//236	354	EC	11101100	ì	&#236;	&igrave;	Latin small letter i with grave
//237	355	ED	11101101	í	&#237;	&iacute;	Latin small letter i with acute
//238	356	EE	11101110	î	&#238;	&icirc;	Latin small letter i with circumflex
//239	357	EF	11101111	ï	&#239;	&iuml;	Latin small letter i with diaeresis
//240	360	F0	11110000	ð	&#240;	&eth;	Latin small letter eth
//241	361	F1	11110001	ñ	&#241;	&ntilde;	Latin small letter n with tilde
//242	362	F2	11110010	ò	&#242;	&ograve;	Latin small letter o with grave
//243	363	F3	11110011	ó	&#243;	&oacute;	Latin small letter o with acute
//244	364	F4	11110100	ô	&#244;	&ocirc;	Latin small letter o with circumflex
//245	365	F5	11110101	õ	&#245;	&otilde;	Latin small letter o with tilde
//246	366	F6	11110110	ö	&#246;	&ouml;	Latin small letter o with diaeresis
//247	367	F7	11110111	÷	&#247;	&divide;	Division sign
//248	370	F8	11111000	ø	&#248;	&oslash;	Latin small letter o with slash
//249	371	F9	11111001	ù	&#249;	&ugrave;	Latin small letter u with grave
//250	372	FA	11111010	ú	&#250;	&uacute;	Latin small letter u with acute
//251	373	FB	11111011	û	&#251;	&ucirc;	Latin small letter u with circumflex
//252	374	FC	11111100	ü	&#252;	&uuml;	Latin small letter u with diaeresis
//253	375	FD	11111101	ý	&#253;	&yacute;	Latin small letter y with acute
//254	376	FE	11111110	þ	&#254;	&thorn;	Latin small letter thorn
//255	377	FF	11111111	ÿ	&#255;	&yuml;	Latin small letter y with diaeresis
